MACRO rom_512x16A
  PIN A[0]
    AntennaGateArea  0.039 ;
  END A[0]
  PIN A[1]
    AntennaGateArea  0.039 ;
  END A[1]
  PIN A[2]
    AntennaGateArea  0.039 ;
  END A[2]
  PIN A[3]
    AntennaGateArea  0.039 ;
  END A[3]
  PIN A[4]
    AntennaGateArea  0.039 ;
  END A[4]
  PIN A[5]
    AntennaGateArea  0.039 ;
  END A[5]
  PIN A[6]
    AntennaGateArea  0.039 ;
  END A[6]
  PIN A[7]
    AntennaGateArea  0.039 ;
  END A[7]
  PIN A[8]
    AntennaGateArea  0.039 ;
  END A[8]
  PIN CEN
    AntennaGateArea  0.039 ;
  END CEN
  PIN CLK
    AntennaGateArea  0.039 ;
  END CLK
END rom_512x16A

END LIBRARY

