
#******
# Preview export LEF
#
#	 Preview sub-version 5.10.41_USR2.19.52
#
# TECH LIB NAME: testLib4
# TECH FILE NAME: techfile.cds
#******

VERSION 5.4 ;

NAMESCASESENSITIVE ON ;

DIVIDERCHAR "|" ;
BUSBITCHARS "<>" ;

 USEMINSPACING OBS OFF  ;
UNITS
    DATABASE MICRONS 2000  ;
END UNITS

 MANUFACTURINGGRID    0.005000 ;

MACRO HEAD8DM
    CLASS CORE ;
    FOREIGN HEAD8DM 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 5.2000 BY 2.8700 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN SLEEP
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.7000 0.7550 2.0150 1.3950 ;
        END
    END SLEEP
    PIN SLEEPOUT
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.1000 0.4950 0.3200 2.4000 ;
        END
    END SLEEPOUT
    PIN VDDG
        DIRECTION INPUT ;
        USE POWER ;
        PORT
        LAYER METAL2 ;
        RECT  2.2000 0.6750 4.5400 1.3950 ;
        END
    END VDDG
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.0000 2.6900 5.2000 3.0500 ;
        RECT  4.8200 1.6700 5.1000 3.0500 ;
        RECT  3.7400 1.6700 4.0200 3.0500 ;
        RECT  2.7000 1.6700 2.9800 3.0500 ;
        RECT  1.6200 2.3950 1.9000 3.0500 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.0000 -0.1800 5.2000 0.1800 ;
        RECT  0.6200 -0.1800 1.3000 0.3200 ;
        RECT  0.6200 -0.1800 0.9000 0.8600 ;
        END
    END VSS
    OBS
        LAYER METAL1 ;
        RECT  4.2600 0.6750 4.5400 2.4300 ;
        RECT  0.6200 2.0400 2.5200 2.2000 ;
        RECT  0.5000 1.1150 1.4600 1.3950 ;
        RECT  1.2200 0.6950 1.4600 1.8550 ;
        RECT  1.1800 1.1150 1.4600 1.8550 ;
        RECT  2.2000 0.6750 2.5200 2.4300 ;
        RECT  2.2000 0.6750 4.5400 1.3950 ;
        RECT  3.2200 0.6750 3.5000 2.4300 ;
        RECT  0.6200 1.6700 0.9000 2.4000 ;
    END
END HEAD8DM

MACRO HEAD16DM
    CLASS CORE ;
    FOREIGN HEAD8DM 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 8.0000 BY 2.8700 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN SLEEP
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.7000 0.7550 2.0150 1.3950 ;
        END
    END SLEEP
    PIN SLEEPOUT
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.1000 0.4950 0.3200 2.4000 ;
        END
    END SLEEPOUT
    PIN VDDG
        DIRECTION INPUT ;
        USE POWER ;
        PORT
        LAYER METAL2 ;
        RECT  2.2000 0.6750 4.5400 1.3950 ;
        END
    END VDDG
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.0000 2.6900 8.0000 3.0500 ;
        RECT  4.7800 1.6700 5.0600 3.0500 ;
        RECT  3.7400 1.6700 4.0200 3.0500 ;
        RECT  2.7000 1.6700 2.9800 3.0500 ;
        RECT  1.6200 2.3950 1.9000 3.0500 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.0000 -0.1800 8.0000 0.1800 ;
        RECT  0.6200 -0.1800 1.3000 0.3200 ;
        RECT  0.6200 -0.1800 0.9000 0.8600 ;
        END
    END VSS
    OBS
        LAYER METAL1 ;
        RECT  7.3800 0.6750 7.6600 2.4300 ;
        RECT  6.3400 0.6750 6.6200 2.4300 ;
        RECT  5.3000 0.6750 5.5800 2.4300 ;
        RECT  4.2600 0.6750 4.5400 2.4300 ;
        RECT  0.6200 2.0400 2.5200 2.2000 ;
        RECT  0.5000 1.1150 1.4600 1.3950 ;
        RECT  1.2200 0.6950 1.4600 1.8550 ;
        RECT  1.1800 1.1150 1.4600 1.8550 ;
        RECT  2.2000 0.6750 2.5200 2.4300 ;
        RECT  2.2000 0.6750 7.6600 1.3950 ;
        RECT  3.2200 0.6750 3.5000 2.4300 ;
        RECT  0.6200 1.6700 0.9000 2.4000 ;
    END
END HEAD16DM

MACRO HEAD32DM
    CLASS CORE ;
    FOREIGN HEAD8DM 0 0 ;
    ORIGIN 0.0000 0.0000 ;
    SIZE 12.0000 BY 2.8700 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN SLEEP
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.7000 0.7550 2.0150 1.3950 ;
        END
    END SLEEP
    PIN SLEEPOUT
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.1000 0.4950 0.3200 2.4000 ;
        END
    END SLEEPOUT
    PIN VDDG
        DIRECTION INPUT ;
        USE POWER ;
        PORT
        LAYER METAL2 ;
        RECT  2.2000 0.6750 4.5400 1.3950 ;
        END
    END VDDG
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.0000 2.6900 12.0000 3.0500 ;
        RECT  4.7800 1.6700 5.0600 3.0500 ;
        RECT  3.7400 1.6700 4.0200 3.0500 ;
        RECT  2.7000 1.6700 2.9800 3.0500 ;
        RECT  1.6200 2.3950 1.9000 3.0500 ;
        END
    END VDD
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.0000 -0.1800 12.0000 0.1800 ;
        RECT  0.6200 -0.1800 1.3000 0.3200 ;
        RECT  0.6200 -0.1800 0.9000 0.8600 ;
        END
    END VSS
    OBS
        LAYER METAL1 ;
        RECT  11.5400 0.6750 11.8200 2.4300 ;
        RECT  10.5000 0.6750 10.7800 2.4300 ;
        RECT  9.4600 0.6750 9.7400 2.4300 ;
        RECT  8.4200 0.6750 8.7000 2.4300 ;
        RECT  7.3800 0.6750 7.6600 2.4300 ;
        RECT  6.3400 0.6750 6.6200 2.4300 ;
        RECT  5.3000 0.6750 5.5800 2.4300 ;
        RECT  4.2600 0.6750 4.5400 2.4300 ;
        RECT  0.6200 2.0400 2.5200 2.2000 ;
        RECT  0.5000 1.1150 1.4600 1.3950 ;
        RECT  1.2200 0.6950 1.4600 1.8550 ;
        RECT  1.1800 1.1150 1.4600 1.8550 ;
        RECT  2.2000 0.6750 2.5200 2.4300 ;
        RECT  2.2000 0.6750 11.6600 1.3950 ;
        RECT  3.2200 0.6750 3.5000 2.4300 ;
        RECT  0.6200 1.6700 0.9000 2.4000 ;
    END
END HEAD32DM

END LIBRARY
