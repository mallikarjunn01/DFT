VERSION 5.4 ;
MACRO ram_256x16A
  PIN A[0]
    ANTENNAGATEAREA  0.039 ;
  END A[0]
  PIN A[1]
    ANTENNAGATEAREA  0.039 ;
  END A[1]
  PIN A[2]
    ANTENNAGATEAREA  0.039 ;
  END A[2]
  PIN A[3]
    ANTENNAGATEAREA  0.039 ;
  END A[3]
  PIN A[4]
    ANTENNAGATEAREA  0.039 ;
  END A[4]
  PIN A[5]
    ANTENNAGATEAREA  0.039 ;
  END A[5]
  PIN A[6]
    ANTENNAGATEAREA  0.039 ;
  END A[6]
  PIN A[7]
    ANTENNAGATEAREA  0.039 ;
  END A[7]
  PIN CEN
    ANTENNAGATEAREA  0.039 ;
  END CEN
  PIN CLK
    ANTENNAGATEAREA  0.039 ;
  END CLK
  PIN D[0]
    ANTENNAGATEAREA  0.039 ;
  END D[0]
  PIN D[10]
    ANTENNAGATEAREA  0.039 ;
  END D[10]
  PIN D[11]
    ANTENNAGATEAREA  0.039 ;
  END D[11]
  PIN D[12]
    ANTENNAGATEAREA  0.039 ;
  END D[12]
  PIN D[13]
    ANTENNAGATEAREA  0.039 ;
  END D[13]
  PIN D[14]
    ANTENNAGATEAREA  0.039 ;
  END D[14]
  PIN D[15]
    ANTENNAGATEAREA  0.039 ;
  END D[15]
  PIN D[1]
    ANTENNAGATEAREA  0.039 ;
  END D[1]
  PIN D[2]
    ANTENNAGATEAREA  0.039 ;
  END D[2]
  PIN D[3]
    ANTENNAGATEAREA  0.039 ;
  END D[3]
  PIN D[4]
    ANTENNAGATEAREA  0.039 ;
  END D[4]
  PIN D[5]
    ANTENNAGATEAREA  0.039 ;
  END D[5]
  PIN D[6]
    ANTENNAGATEAREA  0.039 ;
  END D[6]
  PIN D[7]
    ANTENNAGATEAREA  0.039 ;
  END D[7]
  PIN D[8]
    ANTENNAGATEAREA  0.039 ;
  END D[8]
  PIN D[9]
    ANTENNAGATEAREA  0.039 ;
  END D[9]
  PIN WEN
    ANTENNAGATEAREA  0.039 ;
  END WEN
END ram_256x16A

END LIBRARY
