# Confidential Information of Artisan Components, Inc.
# Use subject to Artisan Components license.
# Copyright (c) 2003 Artisan Components, Inc.

# ACI Version 2002Q3V1

# Bifilator $Revision: 1.161 $
# ADDED ANTENNAEGATEAREA TO LEF


VERSION 5.4 ;


NAMESCASESENSITIVE ON ;

#BUSBITCHARS "[]" ;

# name: ROM-DIFF-HS ROM Generator|TSMC CL013G Process
# version: 2002Q3V1
# comment: 
# configuration:  -instname "rom_512x16A" -words 512 -bits 16 -frequency 166 -ring_width 8 -code_file "rom_512x16A_verilog.rcf" -mux 8 -drive 6 -top_layer met8 -power_type rings -horiz met3 -vert met4 -cust_comment "" -left_bus_delim "[" -right_bus_delim "]" -pwr_gnd_rename "VDD:VDD,GND:VSS" -prefix "" -pin_space 0.0 -name_case upper -check_instname on -diodes on -inside_ring_type GND

# codefile: rom_512x16A_verilog.rcf


MACRO rom_512x16A
  CLASS RING ;
  FOREIGN rom_512x16A 0 0 ;
  ORIGIN 0 0 ;
  SIZE 226.465 BY 184.645 ;
  SYMMETRY X Y R90 ;
  PIN A[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    AntennaGateArea  0.039 ;
    PORT
      LAYER METAL1 ;
      RECT 84.54 21.52 85.2 22.18 ;
      LAYER METAL2 ;
      RECT 84.54 21.52 85.2 22.18 ;
      LAYER METAL3 ;
      RECT 84.54 21.52 85.2 22.18 ;
      LAYER METAL4 ;
      RECT 84.54 21.52 85.2 22.18 ;
      END
    END A[0]
  PIN A[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    AntennaGateArea  0.039 ;
    PORT
      LAYER METAL1 ;
      RECT 80.44 21.52 81.1 22.18 ;
      LAYER METAL2 ;
      RECT 80.44 21.52 81.1 22.18 ;
      LAYER METAL3 ;
      RECT 80.44 21.52 81.1 22.18 ;
      LAYER METAL4 ;
      RECT 80.44 21.52 81.1 22.18 ;
      END
    END A[1]
  PIN A[2]
    DIRECTION INPUT ;
    AntennaGateArea  0.039 ;
    USE SIGNAL ;
    PORT
      LAYER METAL1 ;
      RECT 76.34 21.52 77 22.18 ;
      LAYER METAL2 ;
      RECT 76.34 21.52 77 22.18 ;
      LAYER METAL3 ;
      RECT 76.34 21.52 77 22.18 ;
      LAYER METAL4 ;
      RECT 76.34 21.52 77 22.18 ;
      END
    END A[2]
  PIN A[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    AntennaGateArea  0.039 ;
    PORT
      LAYER METAL1 ;
      RECT 59.94 21.52 60.6 22.18 ;
      LAYER METAL2 ;
      RECT 59.94 21.52 60.6 22.18 ;
      LAYER METAL3 ;
      RECT 59.94 21.52 60.6 22.18 ;
      LAYER METAL4 ;
      RECT 59.94 21.52 60.6 22.18 ;
      END
    END A[3]
  PIN A[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    AntennaGateArea  0.039 ;
    PORT
      LAYER METAL1 ;
      RECT 55.84 21.52 56.5 22.18 ;
      LAYER METAL2 ;
      RECT 55.84 21.52 56.5 22.18 ;
      LAYER METAL3 ;
      RECT 55.84 21.52 56.5 22.18 ;
      LAYER METAL4 ;
      RECT 55.84 21.52 56.5 22.18 ;
      END
    END A[4]
  PIN A[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    AntennaGateArea  0.039 ;
    PORT
      LAYER METAL1 ;
      RECT 51.74 21.52 52.4 22.18 ;
      LAYER METAL2 ;
      RECT 51.74 21.52 52.4 22.18 ;
      LAYER METAL3 ;
      RECT 51.74 21.52 52.4 22.18 ;
      LAYER METAL4 ;
      RECT 51.74 21.52 52.4 22.18 ;
      END
    END A[5]
  PIN A[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    AntennaGateArea  0.039 ;
    PORT
      LAYER METAL1 ;
      RECT 43.54 21.52 44.2 22.18 ;
      LAYER METAL2 ;
      RECT 43.54 21.52 44.2 22.18 ;
      LAYER METAL3 ;
      RECT 43.54 21.52 44.2 22.18 ;
      LAYER METAL4 ;
      RECT 43.54 21.52 44.2 22.18 ;
      END
    END A[6]
  PIN A[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    AntennaGateArea  0.039 ;
    PORT
      LAYER METAL1 ;
      RECT 39.44 21.52 40.1 22.18 ;
      LAYER METAL2 ;
      RECT 39.44 21.52 40.1 22.18 ;
      LAYER METAL3 ;
      RECT 39.44 21.52 40.1 22.18 ;
      LAYER METAL4 ;
      RECT 39.44 21.52 40.1 22.18 ;
      END
    END A[7]
  PIN A[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    AntennaGateArea  0.039 ;
    PORT
      LAYER METAL1 ;
      RECT 35.34 21.52 36 22.18 ;
      LAYER METAL2 ;
      RECT 35.34 21.52 36 22.18 ;
      LAYER METAL3 ;
      RECT 35.34 21.52 36 22.18 ;
      LAYER METAL4 ;
      RECT 35.34 21.52 36 22.18 ;
      END
    END A[8]
  PIN CEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    AntennaGateArea  0.039 ;
    PORT
      LAYER METAL1 ;
      RECT 93.91 17.2 94.57 17.86 ;
      LAYER METAL2 ;
      RECT 93.91 17.2 94.57 17.86 ;
      LAYER METAL3 ;
      RECT 93.91 17.2 94.57 17.86 ;
      LAYER METAL4 ;
      RECT 93.91 17.2 94.57 17.86 ;
      END
    END CEN
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    AntennaGateArea  0.039 ;
    PORT
      LAYER METAL1 ;
      RECT 97.065 17.2 97.725 17.86 ;
      LAYER METAL2 ;
      RECT 97.065 17.2 97.725 17.86 ;
      LAYER METAL3 ;
      RECT 97.065 17.2 97.725 17.86 ;
      LAYER METAL4 ;
      RECT 97.065 17.2 97.725 17.86 ;
      END
    END CLK
  PIN Q[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL1 ;
      RECT 118.055 17.2 118.715 17.86 ;
      LAYER METAL2 ;
      RECT 118.055 17.2 118.715 17.86 ;
      LAYER METAL3 ;
      RECT 118.055 17.2 118.715 17.86 ;
      LAYER METAL4 ;
      RECT 118.055 17.2 118.715 17.86 ;
      END
    END Q[0]
  PIN Q[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL1 ;
      RECT 175.255 17.2 175.915 17.86 ;
      LAYER METAL2 ;
      RECT 175.255 17.2 175.915 17.86 ;
      LAYER METAL3 ;
      RECT 175.255 17.2 175.915 17.86 ;
      LAYER METAL4 ;
      RECT 175.255 17.2 175.915 17.86 ;
      END
    END Q[10]
  PIN Q[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL1 ;
      RECT 180.375 17.2 181.035 17.86 ;
      LAYER METAL2 ;
      RECT 180.375 17.2 181.035 17.86 ;
      LAYER METAL3 ;
      RECT 180.375 17.2 181.035 17.86 ;
      LAYER METAL4 ;
      RECT 180.375 17.2 181.035 17.86 ;
      END
    END Q[11]
  PIN Q[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL1 ;
      RECT 186.695 17.2 187.355 17.86 ;
      LAYER METAL2 ;
      RECT 186.695 17.2 187.355 17.86 ;
      LAYER METAL3 ;
      RECT 186.695 17.2 187.355 17.86 ;
      LAYER METAL4 ;
      RECT 186.695 17.2 187.355 17.86 ;
      END
    END Q[12]
  PIN Q[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL1 ;
      RECT 191.815 17.2 192.475 17.86 ;
      LAYER METAL2 ;
      RECT 191.815 17.2 192.475 17.86 ;
      LAYER METAL3 ;
      RECT 191.815 17.2 192.475 17.86 ;
      LAYER METAL4 ;
      RECT 191.815 17.2 192.475 17.86 ;
      END
    END Q[13]
  PIN Q[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL1 ;
      RECT 198.135 17.2 198.795 17.86 ;
      LAYER METAL2 ;
      RECT 198.135 17.2 198.795 17.86 ;
      LAYER METAL3 ;
      RECT 198.135 17.2 198.795 17.86 ;
      LAYER METAL4 ;
      RECT 198.135 17.2 198.795 17.86 ;
      END
    END Q[14]
  PIN Q[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL1 ;
      RECT 203.255 17.2 203.915 17.86 ;
      LAYER METAL2 ;
      RECT 203.255 17.2 203.915 17.86 ;
      LAYER METAL3 ;
      RECT 203.255 17.2 203.915 17.86 ;
      LAYER METAL4 ;
      RECT 203.255 17.2 203.915 17.86 ;
      END
    END Q[15]
  PIN Q[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL1 ;
      RECT 123.175 17.2 123.835 17.86 ;
      LAYER METAL2 ;
      RECT 123.175 17.2 123.835 17.86 ;
      LAYER METAL3 ;
      RECT 123.175 17.2 123.835 17.86 ;
      LAYER METAL4 ;
      RECT 123.175 17.2 123.835 17.86 ;
      END
    END Q[1]
  PIN Q[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL1 ;
      RECT 129.495 17.2 130.155 17.86 ;
      LAYER METAL2 ;
      RECT 129.495 17.2 130.155 17.86 ;
      LAYER METAL3 ;
      RECT 129.495 17.2 130.155 17.86 ;
      LAYER METAL4 ;
      RECT 129.495 17.2 130.155 17.86 ;
      END
    END Q[2]
  PIN Q[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL1 ;
      RECT 134.615 17.2 135.275 17.86 ;
      LAYER METAL2 ;
      RECT 134.615 17.2 135.275 17.86 ;
      LAYER METAL3 ;
      RECT 134.615 17.2 135.275 17.86 ;
      LAYER METAL4 ;
      RECT 134.615 17.2 135.275 17.86 ;
      END
    END Q[3]
  PIN Q[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL1 ;
      RECT 140.935 17.2 141.595 17.86 ;
      LAYER METAL2 ;
      RECT 140.935 17.2 141.595 17.86 ;
      LAYER METAL3 ;
      RECT 140.935 17.2 141.595 17.86 ;
      LAYER METAL4 ;
      RECT 140.935 17.2 141.595 17.86 ;
      END
    END Q[4]
  PIN Q[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL1 ;
      RECT 146.055 17.2 146.715 17.86 ;
      LAYER METAL2 ;
      RECT 146.055 17.2 146.715 17.86 ;
      LAYER METAL3 ;
      RECT 146.055 17.2 146.715 17.86 ;
      LAYER METAL4 ;
      RECT 146.055 17.2 146.715 17.86 ;
      END
    END Q[5]
  PIN Q[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL1 ;
      RECT 152.375 17.2 153.035 17.86 ;
      LAYER METAL2 ;
      RECT 152.375 17.2 153.035 17.86 ;
      LAYER METAL3 ;
      RECT 152.375 17.2 153.035 17.86 ;
      LAYER METAL4 ;
      RECT 152.375 17.2 153.035 17.86 ;
      END
    END Q[6]
  PIN Q[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL1 ;
      RECT 157.495 17.2 158.155 17.86 ;
      LAYER METAL2 ;
      RECT 157.495 17.2 158.155 17.86 ;
      LAYER METAL3 ;
      RECT 157.495 17.2 158.155 17.86 ;
      LAYER METAL4 ;
      RECT 157.495 17.2 158.155 17.86 ;
      END
    END Q[7]
  PIN Q[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL1 ;
      RECT 163.815 17.2 164.475 17.86 ;
      LAYER METAL2 ;
      RECT 163.815 17.2 164.475 17.86 ;
      LAYER METAL3 ;
      RECT 163.815 17.2 164.475 17.86 ;
      LAYER METAL4 ;
      RECT 163.815 17.2 164.475 17.86 ;
      END
    END Q[8]
  PIN Q[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER METAL1 ;
      RECT 168.935 17.2 169.595 17.86 ;
      LAYER METAL2 ;
      RECT 168.935 17.2 169.595 17.86 ;
      LAYER METAL3 ;
      RECT 168.935 17.2 169.595 17.86 ;
      LAYER METAL4 ;
      RECT 168.935 17.2 169.595 17.86 ;
      END
    END Q[9]
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE RING ;
    PORT
      LAYER METAL3 ;
      RECT 226.465 176.645 0 184.645 ;
      LAYER METAL3 ;
      RECT 0 0 226.465 8 ;
      LAYER METAL4 ;
      RECT 218.465 0 226.465 184.645 ;
      LAYER METAL4 ;
      RECT 0 184.645 8 0 ;
      END
    END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE RING ;
    PORT
      LAYER METAL3 ;
      RECT 217.865 168.045 8.6 176.045 ;
      LAYER METAL3 ;
      RECT 8.6 8.6 217.865 16.6 ;
      LAYER METAL4 ;
      RECT 209.865 8.6 217.865 176.045 ;
      LAYER METAL4 ;
      RECT 8.6 176.045 16.6 8.6 ;
      END
    END VSS
  OBS
    LAYER OVERLAP ;
    POLYGON 17.2 21.52 91.99 21.52 91.99 17.2 209.265 17.2 209.265 167.445
      17.2 167.445 ;
    LAYER VIA12 ;
    POLYGON 17.2 21.52 91.99 21.52 91.99 17.2 209.265 17.2 209.265 167.445
      17.2 167.445 ;
    LAYER VIA23 ;
    POLYGON 17.2 21.52 91.99 21.52 91.99 17.2 209.265 17.2 209.265 167.445
      17.2 167.445 ;
    LAYER VIA34 ;
    POLYGON 17.2 21.52 91.99 21.52 91.99 17.2 209.265 17.2 209.265 167.445
      17.2 167.445 ;
    LAYER VIA45 ;
    POLYGON 17.2 21.52 91.99 21.52 91.99 17.2 209.265 17.2 209.265 167.445
      17.2 167.445 ;
    LAYER METAL1 ;
    POLYGON 17.2 167.445 17.2 21.52 35.16 21.52 35.16 22.36 36.18 22.36
      36.18 21.52 39.26 21.52 39.26 22.36 40.28 22.36 40.28 21.52 43.36 21.52
      43.36 22.36 44.38 22.36 44.38 21.52 51.56 21.52 51.56 22.36 52.58 22.36
      52.58 21.52 55.66 21.52 55.66 22.36 56.68 22.36 56.68 21.52 59.76 21.52
      59.76 22.36 60.78 22.36 60.78 21.52 76.16 21.52 76.16 22.36 77.18 22.36
      77.18 21.52 80.26 21.52 80.26 22.36 81.28 22.36 81.28 21.52 84.36 21.52
      84.36 22.36 85.38 22.36 85.38 21.52 91.99 21.52 91.99 17.2 93.73 17.2
      93.73 18.04 94.75 18.04 94.75 17.2 96.885 17.2 96.885 18.04
      97.905 18.04 97.905 17.2 117.875 17.2 117.875 18.04 118.895 18.04
      118.895 17.2 122.995 17.2 122.995 18.04 124.015 18.04 124.015 17.2
      129.315 17.2 129.315 18.04 130.335 18.04 130.335 17.2 134.435 17.2
      134.435 18.04 135.455 18.04 135.455 17.2 140.755 17.2 140.755 18.04
      141.775 18.04 141.775 17.2 145.875 17.2 145.875 18.04 146.895 18.04
      146.895 17.2 152.195 17.2 152.195 18.04 153.215 18.04 153.215 17.2
      157.315 17.2 157.315 18.04 158.335 18.04 158.335 17.2 163.635 17.2
      163.635 18.04 164.655 18.04 164.655 17.2 168.755 17.2 168.755 18.04
      169.775 18.04 169.775 17.2 175.075 17.2 175.075 18.04 176.095 18.04
      176.095 17.2 180.195 17.2 180.195 18.04 181.215 18.04 181.215 17.2
      186.515 17.2 186.515 18.04 187.535 18.04 187.535 17.2 191.635 17.2
      191.635 18.04 192.655 18.04 192.655 17.2 197.955 17.2 197.955 18.04
      198.975 18.04 198.975 17.2 203.075 17.2 203.075 18.04 204.095 18.04
      204.095 17.2 209.265 17.2 209.265 167.445 ;
    LAYER METAL2 ;
    POLYGON 17.2 167.445 17.2 21.52 35.13 21.52 35.13 22.39 36.21 22.39
      36.21 21.52 39.23 21.52 39.23 22.39 40.31 22.39 40.31 21.52 43.33 21.52
      43.33 22.39 44.41 22.39 44.41 21.52 51.53 21.52 51.53 22.39 52.61 22.39
      52.61 21.52 55.63 21.52 55.63 22.39 56.71 22.39 56.71 21.52 59.73 21.52
      59.73 22.39 60.81 22.39 60.81 21.52 76.13 21.52 76.13 22.39 77.21 22.39
      77.21 21.52 80.23 21.52 80.23 22.39 81.31 22.39 81.31 21.52 84.33 21.52
      84.33 22.39 85.41 22.39 85.41 21.52 91.99 21.52 91.99 17.2 93.7 17.2
      93.7 18.07 94.78 18.07 94.78 17.2 96.855 17.2 96.855 18.07 97.935 18.07
      97.935 17.2 117.845 17.2 117.845 18.07 118.925 18.07 118.925 17.2
      122.965 17.2 122.965 18.07 124.045 18.07 124.045 17.2 129.285 17.2
      129.285 18.07 130.365 18.07 130.365 17.2 134.405 17.2 134.405 18.07
      135.485 18.07 135.485 17.2 140.725 17.2 140.725 18.07 141.805 18.07
      141.805 17.2 145.845 17.2 145.845 18.07 146.925 18.07 146.925 17.2
      152.165 17.2 152.165 18.07 153.245 18.07 153.245 17.2 157.285 17.2
      157.285 18.07 158.365 18.07 158.365 17.2 163.605 17.2 163.605 18.07
      164.685 18.07 164.685 17.2 168.725 17.2 168.725 18.07 169.805 18.07
      169.805 17.2 175.045 17.2 175.045 18.07 176.125 18.07 176.125 17.2
      180.165 17.2 180.165 18.07 181.245 18.07 181.245 17.2 186.485 17.2
      186.485 18.07 187.565 18.07 187.565 17.2 191.605 17.2 191.605 18.07
      192.685 18.07 192.685 17.2 197.925 17.2 197.925 18.07 199.005 18.07
      199.005 17.2 203.045 17.2 203.045 18.07 204.125 18.07 204.125 17.2
      209.265 17.2 209.265 167.445 ;
    LAYER METAL3 ;
    POLYGON 17.2 167.445 17.2 21.52 35.13 21.52 35.13 22.39 36.21 22.39
      36.21 21.52 39.23 21.52 39.23 22.39 40.31 22.39 40.31 21.52 43.33 21.52
      43.33 22.39 44.41 22.39 44.41 21.52 51.53 21.52 51.53 22.39 52.61 22.39
      52.61 21.52 55.63 21.52 55.63 22.39 56.71 22.39 56.71 21.52 59.73 21.52
      59.73 22.39 60.81 22.39 60.81 21.52 76.13 21.52 76.13 22.39 77.21 22.39
      77.21 21.52 80.23 21.52 80.23 22.39 81.31 22.39 81.31 21.52 84.33 21.52
      84.33 22.39 85.41 22.39 85.41 21.52 91.99 21.52 91.99 17.2 93.7 17.2
      93.7 18.07 94.78 18.07 94.78 17.2 96.855 17.2 96.855 18.07 97.935 18.07
      97.935 17.2 117.845 17.2 117.845 18.07 118.925 18.07 118.925 17.2
      122.965 17.2 122.965 18.07 124.045 18.07 124.045 17.2 129.285 17.2
      129.285 18.07 130.365 18.07 130.365 17.2 134.405 17.2 134.405 18.07
      135.485 18.07 135.485 17.2 140.725 17.2 140.725 18.07 141.805 18.07
      141.805 17.2 145.845 17.2 145.845 18.07 146.925 18.07 146.925 17.2
      152.165 17.2 152.165 18.07 153.245 18.07 153.245 17.2 157.285 17.2
      157.285 18.07 158.365 18.07 158.365 17.2 163.605 17.2 163.605 18.07
      164.685 18.07 164.685 17.2 168.725 17.2 168.725 18.07 169.805 18.07
      169.805 17.2 175.045 17.2 175.045 18.07 176.125 18.07 176.125 17.2
      180.165 17.2 180.165 18.07 181.245 18.07 181.245 17.2 186.485 17.2
      186.485 18.07 187.565 18.07 187.565 17.2 191.605 17.2 191.605 18.07
      192.685 18.07 192.685 17.2 197.925 17.2 197.925 18.07 199.005 18.07
      199.005 17.2 203.045 17.2 203.045 18.07 204.125 18.07 204.125 17.2
      209.265 17.2 209.265 167.445 ;
    LAYER METAL4 ;
    POLYGON 17.2 167.445 17.2 21.52 35.13 21.52 35.13 22.39 36.21 22.39
      36.21 21.52 39.23 21.52 39.23 22.39 40.31 22.39 40.31 21.52 43.33 21.52
      43.33 22.39 44.41 22.39 44.41 21.52 51.53 21.52 51.53 22.39 52.61 22.39
      52.61 21.52 55.63 21.52 55.63 22.39 56.71 22.39 56.71 21.52 59.73 21.52
      59.73 22.39 60.81 22.39 60.81 21.52 76.13 21.52 76.13 22.39 77.21 22.39
      77.21 21.52 80.23 21.52 80.23 22.39 81.31 22.39 81.31 21.52 84.33 21.52
      84.33 22.39 85.41 22.39 85.41 21.52 91.99 21.52 91.99 17.2 93.7 17.2
      93.7 18.07 94.78 18.07 94.78 17.2 96.855 17.2 96.855 18.07 97.935 18.07
      97.935 17.2 117.845 17.2 117.845 18.07 118.925 18.07 118.925 17.2
      122.965 17.2 122.965 18.07 124.045 18.07 124.045 17.2 129.285 17.2
      129.285 18.07 130.365 18.07 130.365 17.2 134.405 17.2 134.405 18.07
      135.485 18.07 135.485 17.2 140.725 17.2 140.725 18.07 141.805 18.07
      141.805 17.2 145.845 17.2 145.845 18.07 146.925 18.07 146.925 17.2
      152.165 17.2 152.165 18.07 153.245 18.07 153.245 17.2 157.285 17.2
      157.285 18.07 158.365 18.07 158.365 17.2 163.605 17.2 163.605 18.07
      164.685 18.07 164.685 17.2 168.725 17.2 168.725 18.07 169.805 18.07
      169.805 17.2 175.045 17.2 175.045 18.07 176.125 18.07 176.125 17.2
      180.165 17.2 180.165 18.07 181.245 18.07 181.245 17.2 186.485 17.2
      186.485 18.07 187.565 18.07 187.565 17.2 191.605 17.2 191.605 18.07
      192.685 18.07 192.685 17.2 197.925 17.2 197.925 18.07 199.005 18.07
      199.005 17.2 203.045 17.2 203.045 18.07 204.125 18.07 204.125 17.2
      209.265 17.2 209.265 167.445 ;
    LAYER VIA34 ;
    RECT 209.93 168.11 217.8 175.98 ;
    LAYER VIA34 ;
    RECT 8.665 8.665 16.535 16.535 ;
    LAYER VIA34 ;
    RECT 209.93 8.665 217.8 16.535 ;
    LAYER VIA34 ;
    RECT 8.665 168.11 16.535 175.98 ;
    LAYER VIA34 ;
    RECT 218.53 176.71 226.4 184.58 ;
    LAYER VIA34 ;
    RECT 0.065 0.065 7.935 7.935 ;
    LAYER VIA34 ;
    RECT 218.53 0.065 226.4 7.935 ;
    LAYER VIA34 ;
    RECT 0.065 176.71 7.935 184.58 ;
    LAYER METAL4 ;
    RECT 20.41 167.445 21.99 184.645 ;
    LAYER METAL4 ;
    RECT 24.57 167.445 26.15 184.645 ;
    LAYER METAL4 ;
    RECT 28.27 167.445 30.77 184.645 ;
    LAYER METAL4 ;
    RECT 36.47 167.445 38.97 184.645 ;
    LAYER METAL4 ;
    RECT 44.67 167.445 47.17 184.645 ;
    LAYER METAL4 ;
    RECT 52.87 167.445 55.37 184.645 ;
    LAYER METAL4 ;
    RECT 61.07 167.445 63.57 184.645 ;
    LAYER METAL4 ;
    RECT 69.27 167.445 71.77 184.645 ;
    LAYER METAL4 ;
    RECT 77.47 167.445 79.97 184.645 ;
    LAYER METAL4 ;
    RECT 85.67 167.445 88.17 184.645 ;
    LAYER METAL4 ;
    RECT 90.49 167.445 93.49 184.645 ;
    LAYER METAL4 ;
    RECT 97.63 167.445 100.63 184.645 ;
    LAYER METAL4 ;
    RECT 104.77 167.445 107.77 184.645 ;
    LAYER METAL4 ;
    RECT 110.85 167.445 112.65 184.645 ;
    LAYER METAL4 ;
    RECT 20.41 21.52 21.99 0 ;
    LAYER METAL4 ;
    RECT 24.57 21.52 26.15 0 ;
    LAYER METAL4 ;
    RECT 28.27 21.52 30.77 0 ;
    LAYER METAL4 ;
    RECT 36.47 21.52 38.97 0 ;
    LAYER METAL4 ;
    RECT 44.67 21.52 47.17 0 ;
    LAYER METAL4 ;
    RECT 52.87 21.52 55.37 0 ;
    LAYER METAL4 ;
    RECT 61.07 21.52 63.57 0 ;
    LAYER METAL4 ;
    RECT 69.27 21.52 71.77 0 ;
    LAYER METAL4 ;
    RECT 77.47 21.52 79.97 0 ;
    LAYER METAL4 ;
    RECT 85.67 21.52 88.17 0 ;
    LAYER METAL4 ;
    RECT 91.99 17.2 93.39 0 ;
    LAYER METAL4 ;
    RECT 98.415 17.2 99.815 0 ;
    LAYER METAL4 ;
    RECT 105 17.2 108 0 ;
    LAYER METAL4 ;
    RECT 110.85 17.2 112.65 0 ;
    LAYER METAL4 ;
    RECT 114.935 17.2 115.515 0 ;
    LAYER METAL4 ;
    RECT 117.015 17.2 117.595 0 ;
    LAYER METAL4 ;
    RECT 119.185 17.2 119.765 0 ;
    LAYER METAL4 ;
    RECT 122.125 17.2 122.705 0 ;
    LAYER METAL4 ;
    RECT 124.295 17.2 124.875 0 ;
    LAYER METAL4 ;
    RECT 126.375 17.2 126.955 0 ;
    LAYER METAL4 ;
    RECT 128.455 17.2 129.035 0 ;
    LAYER METAL4 ;
    RECT 130.625 17.2 131.205 0 ;
    LAYER METAL4 ;
    RECT 133.565 17.2 134.145 0 ;
    LAYER METAL4 ;
    RECT 135.735 17.2 136.315 0 ;
    LAYER METAL4 ;
    RECT 137.815 17.2 138.395 0 ;
    LAYER METAL4 ;
    RECT 139.895 17.2 140.475 0 ;
    LAYER METAL4 ;
    RECT 142.065 17.2 142.645 0 ;
    LAYER METAL4 ;
    RECT 145.005 17.2 145.585 0 ;
    LAYER METAL4 ;
    RECT 147.175 17.2 147.755 0 ;
    LAYER METAL4 ;
    RECT 149.255 17.2 149.835 0 ;
    LAYER METAL4 ;
    RECT 151.335 17.2 151.915 0 ;
    LAYER METAL4 ;
    RECT 153.505 17.2 154.085 0 ;
    LAYER METAL4 ;
    RECT 156.445 17.2 157.025 0 ;
    LAYER METAL4 ;
    RECT 158.615 17.2 159.195 0 ;
    LAYER METAL4 ;
    RECT 160.695 17.2 161.275 0 ;
    LAYER METAL4 ;
    RECT 162.775 17.2 163.355 0 ;
    LAYER METAL4 ;
    RECT 164.945 17.2 165.525 0 ;
    LAYER METAL4 ;
    RECT 167.885 17.2 168.465 0 ;
    LAYER METAL4 ;
    RECT 170.055 17.2 170.635 0 ;
    LAYER METAL4 ;
    RECT 172.135 17.2 172.715 0 ;
    LAYER METAL4 ;
    RECT 174.215 17.2 174.795 0 ;
    LAYER METAL4 ;
    RECT 176.385 17.2 176.965 0 ;
    LAYER METAL4 ;
    RECT 179.325 17.2 179.905 0 ;
    LAYER METAL4 ;
    RECT 181.495 17.2 182.075 0 ;
    LAYER METAL4 ;
    RECT 183.575 17.2 184.155 0 ;
    LAYER METAL4 ;
    RECT 185.655 17.2 186.235 0 ;
    LAYER METAL4 ;
    RECT 187.825 17.2 188.405 0 ;
    LAYER METAL4 ;
    RECT 190.765 17.2 191.345 0 ;
    LAYER METAL4 ;
    RECT 192.935 17.2 193.515 0 ;
    LAYER METAL4 ;
    RECT 195.015 17.2 195.595 0 ;
    LAYER METAL4 ;
    RECT 197.095 17.2 197.675 0 ;
    LAYER METAL4 ;
    RECT 199.265 17.2 199.845 0 ;
    LAYER METAL4 ;
    RECT 202.205 17.2 202.785 0 ;
    LAYER METAL4 ;
    RECT 204.375 17.2 204.955 0 ;
    LAYER METAL4 ;
    RECT 206.455 17.2 207.035 0 ;
    LAYER METAL3 ;
    RECT 209.265 21.085 226.465 22.485 ;
    LAYER METAL3 ;
    RECT 209.265 30.355 226.465 31.755 ;
    LAYER METAL3 ;
    RECT 209.265 32.615 226.465 34.015 ;
    LAYER METAL3 ;
    RECT 209.265 35.225 226.465 35.925 ;
    LAYER METAL3 ;
    RECT 209.265 40.26 226.465 42.74 ;
    LAYER METAL3 ;
    RECT 209.265 45.325 226.465 47.925 ;
    LAYER METAL3 ;
    RECT 209.265 50.515 226.465 51.755 ;
    LAYER METAL3 ;
    RECT 209.265 53.445 226.465 54.555 ;
    LAYER METAL3 ;
    RECT 209.265 57.13 226.465 57.83 ;
    LAYER METAL3 ;
    RECT 209.265 66.59 226.465 67.7 ;
    LAYER METAL3 ;
    RECT 209.265 72.31 226.465 74.11 ;
    LAYER METAL3 ;
    RECT 209.265 80.945 226.465 81.645 ;
    LAYER METAL3 ;
    RECT 209.265 84.125 226.465 85.925 ;
    LAYER METAL3 ;
    RECT 209.265 90.535 226.465 91.645 ;
    LAYER METAL3 ;
    RECT 209.265 100.045 226.465 100.745 ;
    LAYER METAL3 ;
    RECT 209.265 102.845 226.465 103.545 ;
    LAYER METAL3 ;
    RECT 209.265 109.675 226.465 112.075 ;
    LAYER METAL3 ;
    RECT 209.265 113.61 226.465 116.01 ;
    LAYER METAL3 ;
    RECT 17.2 24.88 0 25.58 ;
    LAYER METAL3 ;
    RECT 17.2 32.955 0 33.755 ;
    LAYER METAL3 ;
    RECT 17.2 35.055 0 35.755 ;
    LAYER METAL3 ;
    RECT 17.2 40.37 0 41.61 ;
    LAYER METAL3 ;
    RECT 17.2 43.96 0 46.56 ;
    LAYER METAL3 ;
    RECT 17.2 50.515 0 51.755 ;
    LAYER METAL3 ;
    RECT 17.2 53.445 0 54.555 ;
    LAYER METAL3 ;
    RECT 17.2 57.13 0 57.83 ;
    LAYER METAL3 ;
    RECT 17.2 66.59 0 67.7 ;
    LAYER METAL3 ;
    RECT 17.2 72.31 0 74.11 ;
    LAYER METAL3 ;
    RECT 17.2 80.885 0 81.585 ;
    LAYER METAL3 ;
    RECT 17.2 84.125 0 85.925 ;
    LAYER METAL3 ;
    RECT 17.2 90.535 0 91.645 ;
    LAYER METAL3 ;
    RECT 17.2 100.045 0 100.745 ;
    LAYER METAL3 ;
    RECT 17.2 109.675 0 112.075 ;
    LAYER METAL3 ;
    RECT 17.2 113.61 0 116.01 ;
    LAYER METAL3 ;
    RECT 17.2 124.62 0 125.32 ;
    LAYER METAL3 ;
    RECT 17.2 164.35 0 165.05 ;
    LAYER METAL4 ;
    RECT 22.49 167.445 24.07 176.045 ;
    LAYER METAL4 ;
    RECT 26.77 167.445 27.77 176.045 ;
    LAYER METAL4 ;
    RECT 32.37 167.445 34.87 176.045 ;
    LAYER METAL4 ;
    RECT 40.57 167.445 43.07 176.045 ;
    LAYER METAL4 ;
    RECT 48.77 167.445 51.27 176.045 ;
    LAYER METAL4 ;
    RECT 56.97 167.445 59.47 176.045 ;
    LAYER METAL4 ;
    RECT 65.17 167.445 67.67 176.045 ;
    LAYER METAL4 ;
    RECT 73.37 167.445 75.87 176.045 ;
    LAYER METAL4 ;
    RECT 81.57 167.445 84.07 176.045 ;
    LAYER METAL4 ;
    RECT 94.06 167.445 97.06 176.045 ;
    LAYER METAL4 ;
    RECT 101.2 167.445 104.2 176.045 ;
    LAYER METAL4 ;
    RECT 108.29 167.445 110.24 176.045 ;
    LAYER METAL4 ;
    RECT 113.67 167.445 115.07 176.045 ;
    LAYER METAL4 ;
    RECT 115.635 167.445 118.635 176.045 ;
    LAYER METAL4 ;
    RECT 119.755 167.445 121.755 176.045 ;
    LAYER METAL4 ;
    RECT 122.915 167.445 125.915 176.045 ;
    LAYER METAL4 ;
    RECT 127.075 167.445 130.075 176.045 ;
    LAYER METAL4 ;
    RECT 131.195 167.445 133.195 176.045 ;
    LAYER METAL4 ;
    RECT 134.355 167.445 137.355 176.045 ;
    LAYER METAL4 ;
    RECT 138.515 167.445 141.515 176.045 ;
    LAYER METAL4 ;
    RECT 142.635 167.445 144.635 176.045 ;
    LAYER METAL4 ;
    RECT 145.795 167.445 148.795 176.045 ;
    LAYER METAL4 ;
    RECT 149.955 167.445 152.955 176.045 ;
    LAYER METAL4 ;
    RECT 154.075 167.445 156.075 176.045 ;
    LAYER METAL4 ;
    RECT 157.235 167.445 160.235 176.045 ;
    LAYER METAL4 ;
    RECT 161.395 167.445 164.395 176.045 ;
    LAYER METAL4 ;
    RECT 165.515 167.445 167.515 176.045 ;
    LAYER METAL4 ;
    RECT 168.675 167.445 171.675 176.045 ;
    LAYER METAL4 ;
    RECT 172.835 167.445 175.835 176.045 ;
    LAYER METAL4 ;
    RECT 176.955 167.445 178.955 176.045 ;
    LAYER METAL4 ;
    RECT 180.115 167.445 183.115 176.045 ;
    LAYER METAL4 ;
    RECT 184.275 167.445 187.275 176.045 ;
    LAYER METAL4 ;
    RECT 188.395 167.445 190.395 176.045 ;
    LAYER METAL4 ;
    RECT 191.555 167.445 194.555 176.045 ;
    LAYER METAL4 ;
    RECT 195.715 167.445 198.715 176.045 ;
    LAYER METAL4 ;
    RECT 199.835 167.445 201.835 176.045 ;
    LAYER METAL4 ;
    RECT 202.995 167.445 205.995 176.045 ;
    LAYER METAL4 ;
    RECT 207.005 167.445 208.405 176.045 ;
    LAYER METAL4 ;
    RECT 22.49 21.52 24.07 8.6 ;
    LAYER METAL4 ;
    RECT 26.77 21.52 27.77 8.6 ;
    LAYER METAL4 ;
    RECT 32.37 21.52 34.87 8.6 ;
    LAYER METAL4 ;
    RECT 40.57 21.52 43.07 8.6 ;
    LAYER METAL4 ;
    RECT 48.77 21.52 51.27 8.6 ;
    LAYER METAL4 ;
    RECT 56.97 21.52 59.47 8.6 ;
    LAYER METAL4 ;
    RECT 65.17 21.52 67.67 8.6 ;
    LAYER METAL4 ;
    RECT 73.37 21.52 75.87 8.6 ;
    LAYER METAL4 ;
    RECT 81.57 21.52 84.07 8.6 ;
    LAYER METAL4 ;
    RECT 95.11 17.2 96.51 8.6 ;
    LAYER METAL4 ;
    RECT 101.54 17.2 104.54 8.6 ;
    LAYER METAL4 ;
    RECT 108.46 17.2 110.24 8.6 ;
    LAYER METAL4 ;
    RECT 113.205 17.2 114.405 8.6 ;
    LAYER METAL4 ;
    RECT 115.975 17.2 116.555 8.6 ;
    LAYER METAL4 ;
    RECT 120.345 17.2 121.545 8.6 ;
    LAYER METAL4 ;
    RECT 125.335 17.2 125.915 8.6 ;
    LAYER METAL4 ;
    RECT 127.415 17.2 127.995 8.6 ;
    LAYER METAL4 ;
    RECT 131.785 17.2 132.985 8.6 ;
    LAYER METAL4 ;
    RECT 136.775 17.2 137.355 8.6 ;
    LAYER METAL4 ;
    RECT 138.855 17.2 139.435 8.6 ;
    LAYER METAL4 ;
    RECT 143.225 17.2 144.425 8.6 ;
    LAYER METAL4 ;
    RECT 148.215 17.2 148.795 8.6 ;
    LAYER METAL4 ;
    RECT 150.295 17.2 150.875 8.6 ;
    LAYER METAL4 ;
    RECT 154.665 17.2 155.865 8.6 ;
    LAYER METAL4 ;
    RECT 159.655 17.2 160.235 8.6 ;
    LAYER METAL4 ;
    RECT 161.735 17.2 162.315 8.6 ;
    LAYER METAL4 ;
    RECT 166.105 17.2 167.305 8.6 ;
    LAYER METAL4 ;
    RECT 171.095 17.2 171.675 8.6 ;
    LAYER METAL4 ;
    RECT 173.175 17.2 173.755 8.6 ;
    LAYER METAL4 ;
    RECT 177.545 17.2 178.745 8.6 ;
    LAYER METAL4 ;
    RECT 182.535 17.2 183.115 8.6 ;
    LAYER METAL4 ;
    RECT 184.615 17.2 185.195 8.6 ;
    LAYER METAL4 ;
    RECT 188.985 17.2 190.185 8.6 ;
    LAYER METAL4 ;
    RECT 193.975 17.2 194.555 8.6 ;
    LAYER METAL4 ;
    RECT 196.055 17.2 196.635 8.6 ;
    LAYER METAL4 ;
    RECT 200.425 17.2 201.625 8.6 ;
    LAYER METAL4 ;
    RECT 205.415 17.2 205.995 8.6 ;
    LAYER METAL3 ;
    RECT 209.265 18.295 217.865 19.695 ;
    LAYER METAL3 ;
    RECT 209.265 23.685 217.865 25.085 ;
    LAYER METAL3 ;
    RECT 209.265 37.51 217.865 38.75 ;
    LAYER METAL3 ;
    RECT 209.265 48.825 217.865 49.625 ;
    LAYER METAL3 ;
    RECT 209.265 64.3 217.865 65.41 ;
    LAYER METAL3 ;
    RECT 209.265 68.16 217.865 68.86 ;
    LAYER METAL3 ;
    RECT 209.265 77.125 217.865 77.825 ;
    LAYER METAL3 ;
    RECT 209.265 82.105 217.865 83.215 ;
    LAYER METAL3 ;
    RECT 209.265 89.375 217.865 90.075 ;
    LAYER METAL3 ;
    RECT 209.265 92.765 217.865 93.875 ;
    LAYER METAL3 ;
    RECT 209.265 107.695 217.865 109.215 ;
    LAYER METAL3 ;
    RECT 209.265 118.19 217.865 120.19 ;
    LAYER METAL3 ;
    RECT 209.265 122.72 217.865 124.72 ;
    LAYER METAL3 ;
    RECT 209.265 125.22 217.865 127.22 ;
    LAYER METAL3 ;
    RECT 209.265 127.72 217.865 129.72 ;
    LAYER METAL3 ;
    RECT 209.265 130.22 217.865 132.22 ;
    LAYER METAL3 ;
    RECT 209.265 132.72 217.865 134.72 ;
    LAYER METAL3 ;
    RECT 209.265 135.22 217.865 137.22 ;
    LAYER METAL3 ;
    RECT 209.265 137.72 217.865 139.72 ;
    LAYER METAL3 ;
    RECT 209.265 140.22 217.865 142.22 ;
    LAYER METAL3 ;
    RECT 209.265 142.72 217.865 144.72 ;
    LAYER METAL3 ;
    RECT 209.265 145.22 217.865 147.22 ;
    LAYER METAL3 ;
    RECT 209.265 147.72 217.865 149.72 ;
    LAYER METAL3 ;
    RECT 209.265 150.22 217.865 152.22 ;
    LAYER METAL3 ;
    RECT 209.265 152.72 217.865 154.72 ;
    LAYER METAL3 ;
    RECT 209.265 155.22 217.865 157.22 ;
    LAYER METAL3 ;
    RECT 209.265 157.72 217.865 159.72 ;
    LAYER METAL3 ;
    RECT 209.265 160.22 217.865 162.22 ;
    LAYER METAL3 ;
    RECT 209.265 162.7 217.865 165.7 ;
    LAYER METAL3 ;
    RECT 17.2 27.815 8.6 28.615 ;
    LAYER METAL3 ;
    RECT 17.2 30.495 8.6 32.495 ;
    LAYER METAL3 ;
    RECT 17.2 36.215 8.6 37.455 ;
    LAYER METAL3 ;
    RECT 17.2 48.825 8.6 49.625 ;
    LAYER METAL3 ;
    RECT 17.2 64.3 8.6 65.41 ;
    LAYER METAL3 ;
    RECT 17.2 68.2 8.6 68.9 ;
    LAYER METAL3 ;
    RECT 17.2 77.125 8.6 77.825 ;
    LAYER METAL3 ;
    RECT 17.2 82.105 8.6 83.215 ;
    LAYER METAL3 ;
    RECT 17.2 89.335 8.6 90.035 ;
    LAYER METAL3 ;
    RECT 17.2 92.82 8.6 93.82 ;
    LAYER METAL3 ;
    RECT 17.2 107.815 8.6 109.215 ;
    LAYER METAL3 ;
    RECT 17.2 122.12 8.6 122.82 ;
    LAYER METAL3 ;
    RECT 17.2 127.12 8.6 127.82 ;
    LAYER METAL3 ;
    RECT 17.2 129.62 8.6 130.32 ;
    LAYER METAL3 ;
    RECT 17.2 132.12 8.6 132.82 ;
    LAYER METAL3 ;
    RECT 17.2 134.62 8.6 135.32 ;
    LAYER METAL3 ;
    RECT 17.2 137.12 8.6 137.82 ;
    LAYER METAL3 ;
    RECT 17.2 139.62 8.6 140.32 ;
    LAYER METAL3 ;
    RECT 17.2 142.12 8.6 142.82 ;
    LAYER METAL3 ;
    RECT 17.2 144.62 8.6 145.32 ;
    LAYER METAL3 ;
    RECT 17.2 147.12 8.6 147.82 ;
    LAYER METAL3 ;
    RECT 17.2 149.62 8.6 150.32 ;
    LAYER METAL3 ;
    RECT 17.2 152.12 8.6 152.82 ;
    LAYER METAL3 ;
    RECT 17.2 154.62 8.6 155.32 ;
    LAYER METAL3 ;
    RECT 17.2 157.12 8.6 157.82 ;
    LAYER METAL3 ;
    RECT 17.2 159.62 8.6 160.32 ;
    LAYER METAL3 ;
    RECT 17.2 162.12 8.6 162.82 ;
    LAYER VIA34 ;
    RECT 20.625 176.71 21.775 184.58 ;
    LAYER VIA34 ;
    RECT 24.785 176.71 25.935 184.58 ;
    LAYER VIA34 ;
    RECT 28.465 176.71 30.575 184.58 ;
    LAYER VIA34 ;
    RECT 36.665 176.71 38.775 184.58 ;
    LAYER VIA34 ;
    RECT 44.865 176.71 46.975 184.58 ;
    LAYER VIA34 ;
    RECT 53.065 176.71 55.175 184.58 ;
    LAYER VIA34 ;
    RECT 61.265 176.71 63.375 184.58 ;
    LAYER VIA34 ;
    RECT 69.465 176.71 71.575 184.58 ;
    LAYER VIA34 ;
    RECT 77.665 176.71 79.775 184.58 ;
    LAYER VIA34 ;
    RECT 85.865 176.71 87.975 184.58 ;
    LAYER VIA34 ;
    RECT 90.695 176.71 93.285 184.58 ;
    LAYER VIA34 ;
    RECT 97.835 176.71 100.425 184.58 ;
    LAYER VIA34 ;
    RECT 104.975 176.71 107.565 184.58 ;
    LAYER VIA34 ;
    RECT 110.935 176.71 112.565 184.58 ;
    LAYER VIA34 ;
    RECT 20.625 0.065 21.775 7.935 ;
    LAYER VIA34 ;
    RECT 24.785 0.065 25.935 7.935 ;
    LAYER VIA34 ;
    RECT 28.465 0.065 30.575 7.935 ;
    LAYER VIA34 ;
    RECT 36.665 0.065 38.775 7.935 ;
    LAYER VIA34 ;
    RECT 44.865 0.065 46.975 7.935 ;
    LAYER VIA34 ;
    RECT 53.065 0.065 55.175 7.935 ;
    LAYER VIA34 ;
    RECT 61.265 0.065 63.375 7.935 ;
    LAYER VIA34 ;
    RECT 69.465 0.065 71.575 7.935 ;
    LAYER VIA34 ;
    RECT 77.665 0.065 79.775 7.935 ;
    LAYER VIA34 ;
    RECT 85.865 0.065 87.975 7.935 ;
    LAYER VIA34 ;
    RECT 92.115 0.065 93.265 7.935 ;
    LAYER VIA34 ;
    RECT 98.54 0.065 99.69 7.935 ;
    LAYER VIA34 ;
    RECT 105.205 0.065 107.795 7.935 ;
    LAYER VIA34 ;
    RECT 110.935 0.065 112.565 7.935 ;
    LAYER VIA34 ;
    RECT 115.13 0.065 115.32 7.935 ;
    LAYER VIA34 ;
    RECT 117.21 0.065 117.4 7.935 ;
    LAYER VIA34 ;
    RECT 119.38 0.065 119.57 7.935 ;
    LAYER VIA34 ;
    RECT 122.32 0.065 122.51 7.935 ;
    LAYER VIA34 ;
    RECT 124.49 0.065 124.68 7.935 ;
    LAYER VIA34 ;
    RECT 126.57 0.065 126.76 7.935 ;
    LAYER VIA34 ;
    RECT 128.65 0.065 128.84 7.935 ;
    LAYER VIA34 ;
    RECT 130.82 0.065 131.01 7.935 ;
    LAYER VIA34 ;
    RECT 133.76 0.065 133.95 7.935 ;
    LAYER VIA34 ;
    RECT 135.93 0.065 136.12 7.935 ;
    LAYER VIA34 ;
    RECT 138.01 0.065 138.2 7.935 ;
    LAYER VIA34 ;
    RECT 140.09 0.065 140.28 7.935 ;
    LAYER VIA34 ;
    RECT 142.26 0.065 142.45 7.935 ;
    LAYER VIA34 ;
    RECT 145.2 0.065 145.39 7.935 ;
    LAYER VIA34 ;
    RECT 147.37 0.065 147.56 7.935 ;
    LAYER VIA34 ;
    RECT 149.45 0.065 149.64 7.935 ;
    LAYER VIA34 ;
    RECT 151.53 0.065 151.72 7.935 ;
    LAYER VIA34 ;
    RECT 153.7 0.065 153.89 7.935 ;
    LAYER VIA34 ;
    RECT 156.64 0.065 156.83 7.935 ;
    LAYER VIA34 ;
    RECT 158.81 0.065 159 7.935 ;
    LAYER VIA34 ;
    RECT 160.89 0.065 161.08 7.935 ;
    LAYER VIA34 ;
    RECT 162.97 0.065 163.16 7.935 ;
    LAYER VIA34 ;
    RECT 165.14 0.065 165.33 7.935 ;
    LAYER VIA34 ;
    RECT 168.08 0.065 168.27 7.935 ;
    LAYER VIA34 ;
    RECT 170.25 0.065 170.44 7.935 ;
    LAYER VIA34 ;
    RECT 172.33 0.065 172.52 7.935 ;
    LAYER VIA34 ;
    RECT 174.41 0.065 174.6 7.935 ;
    LAYER VIA34 ;
    RECT 176.58 0.065 176.77 7.935 ;
    LAYER VIA34 ;
    RECT 179.52 0.065 179.71 7.935 ;
    LAYER VIA34 ;
    RECT 181.69 0.065 181.88 7.935 ;
    LAYER VIA34 ;
    RECT 183.77 0.065 183.96 7.935 ;
    LAYER VIA34 ;
    RECT 185.85 0.065 186.04 7.935 ;
    LAYER VIA34 ;
    RECT 188.02 0.065 188.21 7.935 ;
    LAYER VIA34 ;
    RECT 190.96 0.065 191.15 7.935 ;
    LAYER VIA34 ;
    RECT 193.13 0.065 193.32 7.935 ;
    LAYER VIA34 ;
    RECT 195.21 0.065 195.4 7.935 ;
    LAYER VIA34 ;
    RECT 197.29 0.065 197.48 7.935 ;
    LAYER VIA34 ;
    RECT 199.46 0.065 199.65 7.935 ;
    LAYER VIA34 ;
    RECT 202.4 0.065 202.59 7.935 ;
    LAYER VIA34 ;
    RECT 204.57 0.065 204.76 7.935 ;
    LAYER VIA34 ;
    RECT 206.65 0.065 206.84 7.935 ;
    LAYER VIA34 ;
    RECT 218.53 21.21 226.4 22.36 ;
    LAYER VIA34 ;
    RECT 218.53 30.48 226.4 31.63 ;
    LAYER VIA34 ;
    RECT 218.53 32.74 226.4 33.89 ;
    LAYER VIA34 ;
    RECT 218.53 35.48 226.4 35.67 ;
    LAYER VIA34 ;
    RECT 218.53 40.445 226.4 42.555 ;
    LAYER VIA34 ;
    RECT 218.53 45.57 226.4 47.68 ;
    LAYER VIA34 ;
    RECT 218.53 50.8 226.4 51.47 ;
    LAYER VIA34 ;
    RECT 218.53 53.665 226.4 54.335 ;
    LAYER VIA34 ;
    RECT 218.53 57.385 226.4 57.575 ;
    LAYER VIA34 ;
    RECT 218.53 66.81 226.4 67.48 ;
    LAYER VIA34 ;
    RECT 218.53 72.395 226.4 74.025 ;
    LAYER VIA34 ;
    RECT 218.53 81.2 226.4 81.39 ;
    LAYER VIA34 ;
    RECT 218.53 84.21 226.4 85.84 ;
    LAYER VIA34 ;
    RECT 218.53 90.755 226.4 91.425 ;
    LAYER VIA34 ;
    RECT 218.53 100.3 226.4 100.49 ;
    LAYER VIA34 ;
    RECT 218.53 103.1 226.4 103.29 ;
    LAYER VIA34 ;
    RECT 218.53 109.82 226.4 111.93 ;
    LAYER VIA34 ;
    RECT 218.53 113.755 226.4 115.865 ;
    LAYER VIA34 ;
    RECT 0.065 25.135 7.935 25.325 ;
    LAYER VIA34 ;
    RECT 0.065 33.02 7.935 33.69 ;
    LAYER VIA34 ;
    RECT 0.065 35.31 7.935 35.5 ;
    LAYER VIA34 ;
    RECT 0.065 40.655 7.935 41.325 ;
    LAYER VIA34 ;
    RECT 0.065 44.205 7.935 46.315 ;
    LAYER VIA34 ;
    RECT 0.065 50.8 7.935 51.47 ;
    LAYER VIA34 ;
    RECT 0.065 53.665 7.935 54.335 ;
    LAYER VIA34 ;
    RECT 0.065 57.385 7.935 57.575 ;
    LAYER VIA34 ;
    RECT 0.065 66.81 7.935 67.48 ;
    LAYER VIA34 ;
    RECT 0.065 72.395 7.935 74.025 ;
    LAYER VIA34 ;
    RECT 0.065 81.14 7.935 81.33 ;
    LAYER VIA34 ;
    RECT 0.065 84.21 7.935 85.84 ;
    LAYER VIA34 ;
    RECT 0.065 90.755 7.935 91.425 ;
    LAYER VIA34 ;
    RECT 0.065 100.3 7.935 100.49 ;
    LAYER VIA34 ;
    RECT 0.065 109.82 7.935 111.93 ;
    LAYER VIA34 ;
    RECT 0.065 113.755 7.935 115.865 ;
    LAYER VIA34 ;
    RECT 0.065 124.875 7.935 125.065 ;
    LAYER VIA34 ;
    RECT 0.065 164.605 7.935 164.795 ;
    LAYER VIA34 ;
    RECT 22.705 168.11 23.855 175.98 ;
    LAYER VIA34 ;
    RECT 26.935 168.11 27.605 175.98 ;
    LAYER VIA34 ;
    RECT 32.565 168.11 34.675 175.98 ;
    LAYER VIA34 ;
    RECT 40.765 168.11 42.875 175.98 ;
    LAYER VIA34 ;
    RECT 48.965 168.11 51.075 175.98 ;
    LAYER VIA34 ;
    RECT 57.165 168.11 59.275 175.98 ;
    LAYER VIA34 ;
    RECT 65.365 168.11 67.475 175.98 ;
    LAYER VIA34 ;
    RECT 73.565 168.11 75.675 175.98 ;
    LAYER VIA34 ;
    RECT 81.765 168.11 83.875 175.98 ;
    LAYER VIA34 ;
    RECT 94.265 168.11 96.855 175.98 ;
    LAYER VIA34 ;
    RECT 101.405 168.11 103.995 175.98 ;
    LAYER VIA34 ;
    RECT 108.45 168.11 110.08 175.98 ;
    LAYER VIA34 ;
    RECT 113.795 168.11 114.945 175.98 ;
    LAYER VIA34 ;
    RECT 115.84 168.11 118.43 175.98 ;
    LAYER VIA34 ;
    RECT 119.94 168.11 121.57 175.98 ;
    LAYER VIA34 ;
    RECT 123.12 168.11 125.71 175.98 ;
    LAYER VIA34 ;
    RECT 127.28 168.11 129.87 175.98 ;
    LAYER VIA34 ;
    RECT 131.38 168.11 133.01 175.98 ;
    LAYER VIA34 ;
    RECT 134.56 168.11 137.15 175.98 ;
    LAYER VIA34 ;
    RECT 138.72 168.11 141.31 175.98 ;
    LAYER VIA34 ;
    RECT 142.82 168.11 144.45 175.98 ;
    LAYER VIA34 ;
    RECT 146 168.11 148.59 175.98 ;
    LAYER VIA34 ;
    RECT 150.16 168.11 152.75 175.98 ;
    LAYER VIA34 ;
    RECT 154.26 168.11 155.89 175.98 ;
    LAYER VIA34 ;
    RECT 157.44 168.11 160.03 175.98 ;
    LAYER VIA34 ;
    RECT 161.6 168.11 164.19 175.98 ;
    LAYER VIA34 ;
    RECT 165.7 168.11 167.33 175.98 ;
    LAYER VIA34 ;
    RECT 168.88 168.11 171.47 175.98 ;
    LAYER VIA34 ;
    RECT 173.04 168.11 175.63 175.98 ;
    LAYER VIA34 ;
    RECT 177.14 168.11 178.77 175.98 ;
    LAYER VIA34 ;
    RECT 180.32 168.11 182.91 175.98 ;
    LAYER VIA34 ;
    RECT 184.48 168.11 187.07 175.98 ;
    LAYER VIA34 ;
    RECT 188.58 168.11 190.21 175.98 ;
    LAYER VIA34 ;
    RECT 191.76 168.11 194.35 175.98 ;
    LAYER VIA34 ;
    RECT 195.92 168.11 198.51 175.98 ;
    LAYER VIA34 ;
    RECT 200.02 168.11 201.65 175.98 ;
    LAYER VIA34 ;
    RECT 203.2 168.11 205.79 175.98 ;
    LAYER VIA34 ;
    RECT 207.13 168.11 208.28 175.98 ;
    LAYER VIA34 ;
    RECT 22.705 8.665 23.855 16.535 ;
    LAYER VIA34 ;
    RECT 26.935 8.665 27.605 16.535 ;
    LAYER VIA34 ;
    RECT 32.565 8.665 34.675 16.535 ;
    LAYER VIA34 ;
    RECT 40.765 8.665 42.875 16.535 ;
    LAYER VIA34 ;
    RECT 48.965 8.665 51.075 16.535 ;
    LAYER VIA34 ;
    RECT 57.165 8.665 59.275 16.535 ;
    LAYER VIA34 ;
    RECT 65.365 8.665 67.475 16.535 ;
    LAYER VIA34 ;
    RECT 73.565 8.665 75.675 16.535 ;
    LAYER VIA34 ;
    RECT 81.765 8.665 83.875 16.535 ;
    LAYER VIA34 ;
    RECT 95.235 8.665 96.385 16.535 ;
    LAYER VIA34 ;
    RECT 101.745 8.665 104.335 16.535 ;
    LAYER VIA34 ;
    RECT 108.535 8.665 110.165 16.535 ;
    LAYER VIA34 ;
    RECT 113.47 8.665 114.14 16.535 ;
    LAYER VIA34 ;
    RECT 116.17 8.665 116.36 16.535 ;
    LAYER VIA34 ;
    RECT 120.61 8.665 121.28 16.535 ;
    LAYER VIA34 ;
    RECT 125.53 8.665 125.72 16.535 ;
    LAYER VIA34 ;
    RECT 127.61 8.665 127.8 16.535 ;
    LAYER VIA34 ;
    RECT 132.05 8.665 132.72 16.535 ;
    LAYER VIA34 ;
    RECT 136.97 8.665 137.16 16.535 ;
    LAYER VIA34 ;
    RECT 139.05 8.665 139.24 16.535 ;
    LAYER VIA34 ;
    RECT 143.49 8.665 144.16 16.535 ;
    LAYER VIA34 ;
    RECT 148.41 8.665 148.6 16.535 ;
    LAYER VIA34 ;
    RECT 150.49 8.665 150.68 16.535 ;
    LAYER VIA34 ;
    RECT 154.93 8.665 155.6 16.535 ;
    LAYER VIA34 ;
    RECT 159.85 8.665 160.04 16.535 ;
    LAYER VIA34 ;
    RECT 161.93 8.665 162.12 16.535 ;
    LAYER VIA34 ;
    RECT 166.37 8.665 167.04 16.535 ;
    LAYER VIA34 ;
    RECT 171.29 8.665 171.48 16.535 ;
    LAYER VIA34 ;
    RECT 173.37 8.665 173.56 16.535 ;
    LAYER VIA34 ;
    RECT 177.81 8.665 178.48 16.535 ;
    LAYER VIA34 ;
    RECT 182.73 8.665 182.92 16.535 ;
    LAYER VIA34 ;
    RECT 184.81 8.665 185 16.535 ;
    LAYER VIA34 ;
    RECT 189.25 8.665 189.92 16.535 ;
    LAYER VIA34 ;
    RECT 194.17 8.665 194.36 16.535 ;
    LAYER VIA34 ;
    RECT 196.25 8.665 196.44 16.535 ;
    LAYER VIA34 ;
    RECT 200.69 8.665 201.36 16.535 ;
    LAYER VIA34 ;
    RECT 205.61 8.665 205.8 16.535 ;
    LAYER VIA34 ;
    RECT 209.93 18.42 217.8 19.57 ;
    LAYER VIA34 ;
    RECT 209.93 23.81 217.8 24.96 ;
    LAYER VIA34 ;
    RECT 209.93 37.795 217.8 38.465 ;
    LAYER VIA34 ;
    RECT 209.93 48.89 217.8 49.56 ;
    LAYER VIA34 ;
    RECT 209.93 64.52 217.8 65.19 ;
    LAYER VIA34 ;
    RECT 209.93 68.415 217.8 68.605 ;
    LAYER VIA34 ;
    RECT 209.93 77.38 217.8 77.57 ;
    LAYER VIA34 ;
    RECT 209.93 82.325 217.8 82.995 ;
    LAYER VIA34 ;
    RECT 209.93 89.63 217.8 89.82 ;
    LAYER VIA34 ;
    RECT 209.93 92.985 217.8 93.655 ;
    LAYER VIA34 ;
    RECT 209.93 107.88 217.8 109.03 ;
    LAYER VIA34 ;
    RECT 209.93 118.375 217.8 120.005 ;
    LAYER VIA34 ;
    RECT 209.93 122.905 217.8 124.535 ;
    LAYER VIA34 ;
    RECT 209.93 125.405 217.8 127.035 ;
    LAYER VIA34 ;
    RECT 209.93 127.905 217.8 129.535 ;
    LAYER VIA34 ;
    RECT 209.93 130.405 217.8 132.035 ;
    LAYER VIA34 ;
    RECT 209.93 132.905 217.8 134.535 ;
    LAYER VIA34 ;
    RECT 209.93 135.405 217.8 137.035 ;
    LAYER VIA34 ;
    RECT 209.93 137.905 217.8 139.535 ;
    LAYER VIA34 ;
    RECT 209.93 140.405 217.8 142.035 ;
    LAYER VIA34 ;
    RECT 209.93 142.905 217.8 144.535 ;
    LAYER VIA34 ;
    RECT 209.93 145.405 217.8 147.035 ;
    LAYER VIA34 ;
    RECT 209.93 147.905 217.8 149.535 ;
    LAYER VIA34 ;
    RECT 209.93 150.405 217.8 152.035 ;
    LAYER VIA34 ;
    RECT 209.93 152.905 217.8 154.535 ;
    LAYER VIA34 ;
    RECT 209.93 155.405 217.8 157.035 ;
    LAYER VIA34 ;
    RECT 209.93 157.905 217.8 159.535 ;
    LAYER VIA34 ;
    RECT 209.93 160.405 217.8 162.035 ;
    LAYER VIA34 ;
    RECT 209.93 162.905 217.8 165.495 ;
    LAYER VIA34 ;
    RECT 8.665 27.88 16.535 28.55 ;
    LAYER VIA34 ;
    RECT 8.665 30.68 16.535 32.31 ;
    LAYER VIA34 ;
    RECT 8.665 36.5 16.535 37.17 ;
    LAYER VIA34 ;
    RECT 8.665 48.89 16.535 49.56 ;
    LAYER VIA34 ;
    RECT 8.665 64.52 16.535 65.19 ;
    LAYER VIA34 ;
    RECT 8.665 68.455 16.535 68.645 ;
    LAYER VIA34 ;
    RECT 8.665 77.38 16.535 77.57 ;
    LAYER VIA34 ;
    RECT 8.665 82.325 16.535 82.995 ;
    LAYER VIA34 ;
    RECT 8.665 89.59 16.535 89.78 ;
    LAYER VIA34 ;
    RECT 8.665 92.985 16.535 93.655 ;
    LAYER VIA34 ;
    RECT 8.665 107.94 16.535 109.09 ;
    LAYER VIA34 ;
    RECT 8.665 122.375 16.535 122.565 ;
    LAYER VIA34 ;
    RECT 8.665 127.375 16.535 127.565 ;
    LAYER VIA34 ;
    RECT 8.665 129.875 16.535 130.065 ;
    LAYER VIA34 ;
    RECT 8.665 132.375 16.535 132.565 ;
    LAYER VIA34 ;
    RECT 8.665 134.875 16.535 135.065 ;
    LAYER VIA34 ;
    RECT 8.665 137.375 16.535 137.565 ;
    LAYER VIA34 ;
    RECT 8.665 139.875 16.535 140.065 ;
    LAYER VIA34 ;
    RECT 8.665 142.375 16.535 142.565 ;
    LAYER VIA34 ;
    RECT 8.665 144.875 16.535 145.065 ;
    LAYER VIA34 ;
    RECT 8.665 147.375 16.535 147.565 ;
    LAYER VIA34 ;
    RECT 8.665 149.875 16.535 150.065 ;
    LAYER VIA34 ;
    RECT 8.665 152.375 16.535 152.565 ;
    LAYER VIA34 ;
    RECT 8.665 154.875 16.535 155.065 ;
    LAYER VIA34 ;
    RECT 8.665 157.375 16.535 157.565 ;
    LAYER VIA34 ;
    RECT 8.665 159.875 16.535 160.065 ;
    LAYER VIA34 ;
    RECT 8.665 162.375 16.535 162.565 ;
    END
  #BEGINEXT "VSI SIGNATURE 1.0"
    #CREATOR "Artisan Components, Inc." ;
    #DATE "2003-10-27" ;
    #REVISION "1.0" ;
    #ENDEXT
  END rom_512x16A
END LIBRARY

