#----------------------------------------------------------------------------
# Copyright (C) 2002 Taiwan Semiconductor Manufacturing Company, Ltd.
# Confidential Information of TSMC, Ltd.
# Use subject to TSMC Design Service Division license.
#
# Input source : ANTENNA.DB
# File         : antenna.lef
# Date         : Tue Jul 16 21:08:53 2002
#----------------------------------------------------------------------------
# TSMC Antenna Rule for Silicon Ensemble v5.3
#----------------------------------------------------------------------------
#
#     "AntennaGateArea" is derived from W, L parameters of MOS transistor. 
#  Since Silicon Ensemble v5.3 is improved to know diffusion diode area,
#  AD/AS and diode area parameter will be used for "AntennaDiffArea". 
#
#    Notice that this antenna rule only works for Silicon Ensemble v5.3 and
#  after. For detail information, please refer to Cadence application note -
# "Detail Calculation of Process Antenna Effect".
#
#-----------------------------------------------------------------------------

LAYER METAL1
    Thickness 0.260000 ;
    AntennaCumAreaRatio 600.000000 ;
    AntennaCumDiffAreaRatio PWL ( ( 0 600 ) ( 0.159 600 ) ( 0.160 43072.96 ) ( 0.5 43228 ) ( 1 43456 ) ( 1.5 43684 ) ) ;
END METAL1

LAYER METAL2
    Thickness 0.350000 ;
    AntennaCumAreaRatio 600.000000 ;
    AntennaCumDiffAreaRatio PWL ( ( 0 600 ) ( 0.159 600 ) ( 0.160 43072.96 ) ( 0.5 43228 ) ( 1 43456 ) ( 1.5 43684 ) ) ;
END METAL2

LAYER METAL3
    Thickness 0.350000 ;
    AntennaCumAreaRatio 600.000000 ;
    AntennaCumDiffAreaRatio PWL ( ( 0 600 ) ( 0.159 600 ) ( 0.160 43072.96 ) ( 0.5 43228 ) ( 1 43456 ) ( 1.5 43684 ) ) ;
END METAL3

LAYER METAL4
    Thickness 0.350000 ;
    AntennaCumAreaRatio 600.000000 ;
    AntennaCumDiffAreaRatio PWL ( ( 0 600 ) ( 0.159 600 ) ( 0.160 43072.96 ) ( 0.5 43228 ) ( 1 43456 ) ( 1.5 43684 ) ) ;
END METAL4

LAYER METAL5
    Thickness 0.350000 ;
    AntennaCumAreaRatio 600.000000 ;
    AntennaCumDiffAreaRatio PWL ( ( 0 600 ) ( 0.159 600 ) ( 0.160 43072.96 ) ( 0.5 43228 ) ( 1 43456 ) ( 1.5 43684 ) ) ;
END METAL5

LAYER METAL6
    Thickness 0.350000 ;
    AntennaCumAreaRatio 600.000000 ;
    AntennaCumDiffAreaRatio PWL ( ( 0 600 ) ( 0.159 600 ) ( 0.160 43072.96 ) ( 0.5 43228 ) ( 1 43456 ) ( 1.5 43684 ) ) ;
END METAL6

LAYER METAL7
    Thickness 0.900000 ;
    AntennaCumAreaRatio 600.000000 ;
    AntennaCumDiffAreaRatio PWL ( ( 0 600 ) ( 0.159 600 ) ( 0.160 51280 ) ( 0.5 54000 ) ( 1 58000 ) ( 1.5 62000 ) ) ;
END METAL7

LAYER VIA12
    AntennaAreaRatio 20.000000 ;
    AntennaDiffAreaRatio PWL ( ( 0 20 ) ( 0.159 20 ) (0.160 933.6 ) ( 0.5 1005 ) ( 1 1110 ) ( 1.5 1215 ) ) ;
END VIA12

LAYER VIA23
    AntennaAreaRatio 20.000000 ;
    AntennaDiffAreaRatio PWL ( ( 0 20 ) ( 0.159 20 ) (0.160 933.6 ) ( 0.5 1005 ) ( 1 1110 ) ( 1.5 1215 ) ) ;
END VIA23

LAYER VIA34
    AntennaAreaRatio 20.000000 ;
    AntennaDiffAreaRatio PWL ( ( 0 20 ) ( 0.159 20 ) (0.160 933.6 ) ( 0.5 1005 ) ( 1 1110 ) ( 1.5 1215 ) ) ;
END VIA34

LAYER VIA45
    AntennaAreaRatio 20.000000 ;
    AntennaDiffAreaRatio PWL ( ( 0 20 ) ( 0.159 20 ) (0.160 933.6 ) ( 0.5 1005 ) ( 1 1110 ) ( 1.5 1215 ) ) ;
END VIA45

LAYER VIA56
    AntennaAreaRatio 20.000000 ;
    AntennaDiffAreaRatio PWL ( ( 0 20 ) ( 0.159 20 ) (0.160 933.6 ) ( 0.5 1005 ) ( 1 1110 ) ( 1.5 1215 ) ) ;
END VIA56

LAYER VIA67
    AntennaAreaRatio 20.000000 ;
    AntennaDiffAreaRatio PWL ( ( 0 20 ) ( 0.159 20 ) (0.160 933.6 ) ( 0.5 1005 ) ( 1 1110 ) ( 1.5 1215 ) ) ;
END VIA67

MACRO PDD12DGZ
    PIN C
        AntennaDiffArea 3.660000 ;
    END C
    PIN I
        AntennaGateArea 2.600000 ;
    END I
    PIN OEN
        AntennaGateArea 2.730000 ;
    END OEN
    PIN PAD
        AntennaGateArea 3.600000 ;
        AntennaDiffArea 3478.000000 ;
    END PAD
END PDD12DGZ

MACRO PDUSDGZ
    PIN C
        AntennaDiffArea 3.660000 ;
    END C
    PIN PAD
        AntennaGateArea 4.800000 ;
        AntennaDiffArea 3670.000000 ;
    END PAD
END PDUSDGZ

MACRO PDB24DGZ
    PIN C
        AntennaDiffArea 3.660000 ;
    END C
    PIN I
        AntennaGateArea 2.600000 ;
    END I
    PIN OEN
        AntennaGateArea 2.730000 ;
    END OEN
    PIN PAD
        AntennaGateArea 3.600000 ;
        AntennaDiffArea 3479.000000 ;
    END PAD
END PDB24DGZ

MACRO PRU24DGZ
    PIN C
        AntennaDiffArea 3.660000 ;
    END C
    PIN I
        AntennaGateArea 2.600000 ;
    END I
    PIN OEN
        AntennaGateArea 2.730000 ;
    END OEN
    PIN PAD
        AntennaGateArea 3.600000 ;
        AntennaDiffArea 3479.000000 ;
    END PAD
END PRU24DGZ

MACRO PDB08DGZ
    PIN C
        AntennaDiffArea 3.660000 ;
    END C
    PIN I
        AntennaGateArea 2.600000 ;
    END I
    PIN OEN
        AntennaGateArea 2.730000 ;
    END OEN
    PIN PAD
        AntennaGateArea 3.600000 ;
        AntennaDiffArea 3486.000000 ;
    END PAD
END PDB08DGZ

MACRO PRU08DGZ
    PIN C
        AntennaDiffArea 3.660000 ;
    END C
    PIN I
        AntennaGateArea 2.600000 ;
    END I
    PIN OEN
        AntennaGateArea 2.730000 ;
    END OEN
    PIN PAD
        AntennaGateArea 3.600000 ;
        AntennaDiffArea 3486.000000 ;
    END PAD
END PRU08DGZ

MACRO PDD16DGZ
    PIN C
        AntennaDiffArea 3.660000 ;
    END C
    PIN I
        AntennaGateArea 2.600000 ;
    END I
    PIN OEN
        AntennaGateArea 2.730000 ;
    END OEN
    PIN PAD
        AntennaGateArea 3.600000 ;
        AntennaDiffArea 3217.000000 ;
    END PAD
END PDD16DGZ

MACRO PRO24CDG
    PIN I
        AntennaGateArea 2.600000 ;
    END I
    PIN PAD
        AntennaDiffArea 4047.000000 ;
    END PAD
END PRO24CDG

MACRO PDUWDGZ
    PIN C
        AntennaDiffArea 3.660000 ;
    END C
    PIN PAD
        AntennaGateArea 3.600000 ;
        AntennaDiffArea 3670.000000 ;
    END PAD
    PIN REN
        AntennaGateArea 8.170000 ;
    END REN
END PDUWDGZ

MACRO PRO08CDG
    PIN I
        AntennaGateArea 2.600000 ;
    END I
    PIN PAD
        AntennaDiffArea 4037.000000 ;
    END PAD
END PRO08CDG

MACRO PRD12DGZ
    PIN C
        AntennaDiffArea 3.660000 ;
    END C
    PIN I
        AntennaGateArea 2.600000 ;
    END I
    PIN OEN
        AntennaGateArea 2.730000 ;
    END OEN
    PIN PAD
        AntennaGateArea 3.600000 ;
        AntennaDiffArea 3478.000000 ;
    END PAD
END PRD12DGZ

MACRO PRB24DGZ
    PIN C
        AntennaDiffArea 3.660000 ;
    END C
    PIN I
        AntennaGateArea 2.600000 ;
    END I
    PIN OEN
        AntennaGateArea 2.730000 ;
    END OEN
    PIN PAD
        AntennaGateArea 3.600000 ;
        AntennaDiffArea 3479.000000 ;
    END PAD
END PRB24DGZ

MACRO PDT02DGZ
    PIN I
        AntennaGateArea 2.600000 ;
    END I
    PIN OEN
        AntennaGateArea 2.730000 ;
    END OEN
    PIN PAD
        AntennaDiffArea 3652.000000 ;
    END PAD
END PDT02DGZ

MACRO PDT12DGZ
    PIN I
        AntennaGateArea 2.600000 ;
    END I
    PIN OEN
        AntennaGateArea 2.730000 ;
    END OEN
    PIN PAD
        AntennaDiffArea 3461.000000 ;
    END PAD
END PDT12DGZ

MACRO PRB08DGZ
    PIN C
        AntennaDiffArea 3.660000 ;
    END C
    PIN I
        AntennaGateArea 2.600000 ;
    END I
    PIN OEN
        AntennaGateArea 2.730000 ;
    END OEN
    PIN PAD
        AntennaGateArea 3.600000 ;
        AntennaDiffArea 3486.000000 ;
    END PAD
END PRB08DGZ

MACRO PRU12SDGZ
    PIN C
        AntennaDiffArea 3.660000 ;
    END C
    PIN I
        AntennaGateArea 2.600000 ;
    END I
    PIN OEN
        AntennaGateArea 2.730000 ;
    END OEN
    PIN PAD
        AntennaGateArea 4.800000 ;
        AntennaDiffArea 3478.000000 ;
    END PAD
END PRU12SDGZ

MACRO PRD16DGZ
    PIN C
        AntennaDiffArea 3.660000 ;
    END C
    PIN I
        AntennaGateArea 2.600000 ;
    END I
    PIN OEN
        AntennaGateArea 2.730000 ;
    END OEN
    PIN PAD
        AntennaGateArea 3.600000 ;
        AntennaDiffArea 3217.000000 ;
    END PAD
END PRD16DGZ

MACRO PDT16DGZ
    PIN I
        AntennaGateArea 2.600000 ;
    END I
    PIN OEN
        AntennaGateArea 2.730000 ;
    END OEN
    PIN PAD
        AntennaDiffArea 3200.000000 ;
    END PAD
END PDT16DGZ

MACRO PDB24SDGZ
    PIN C
        AntennaDiffArea 3.660000 ;
    END C
    PIN I
        AntennaGateArea 2.600000 ;
    END I
    PIN OEN
        AntennaGateArea 2.730000 ;
    END OEN
    PIN PAD
        AntennaGateArea 4.800000 ;
        AntennaDiffArea 3479.000000 ;
    END PAD
END PDB24SDGZ

MACRO PRU16SDGZ
    PIN C
        AntennaDiffArea 3.660000 ;
    END C
    PIN I
        AntennaGateArea 2.600000 ;
    END I
    PIN OEN
        AntennaGateArea 2.730000 ;
    END OEN
    PIN PAD
        AntennaGateArea 4.800000 ;
        AntennaDiffArea 3217.000000 ;
    END PAD
END PRU16SDGZ

MACRO PDD24SDGZ
    PIN C
        AntennaDiffArea 3.660000 ;
    END C
    PIN I
        AntennaGateArea 2.600000 ;
    END I
    PIN OEN
        AntennaGateArea 2.730000 ;
    END OEN
    PIN PAD
        AntennaGateArea 4.800000 ;
        AntennaDiffArea 3479.000000 ;
    END PAD
END PDD24SDGZ

MACRO PDDW04DGZ
    PIN C
        AntennaDiffArea 3.660000 ;
    END C
    PIN I
        AntennaGateArea 2.600000 ;
    END I
    PIN OEN
        AntennaGateArea 2.730000 ;
    END OEN
    PIN PAD
        AntennaGateArea 3.600000 ;
        AntennaDiffArea 3484.000000 ;
    END PAD
    PIN REN
        AntennaGateArea 1.170000 ;
    END REN
END PDDW04DGZ

MACRO PDDW24DGZ
    PIN C
        AntennaDiffArea 3.660000 ;
    END C
    PIN I
        AntennaGateArea 2.600000 ;
    END I
    PIN OEN
        AntennaGateArea 2.730000 ;
    END OEN
    PIN PAD
        AntennaGateArea 3.600000 ;
        AntennaDiffArea 3479.000000 ;
    END PAD
    PIN REN
        AntennaGateArea 1.170000 ;
    END REN
END PDDW24DGZ

MACRO PDDW08DGZ
    PIN C
        AntennaDiffArea 3.660000 ;
    END C
    PIN I
        AntennaGateArea 2.600000 ;
    END I
    PIN OEN
        AntennaGateArea 2.730000 ;
    END OEN
    PIN PAD
        AntennaGateArea 3.600000 ;
        AntennaDiffArea 3486.000000 ;
    END PAD
    PIN REN
        AntennaGateArea 1.170000 ;
    END REN
END PDDW08DGZ

MACRO PRT12DGZ
    PIN I
        AntennaGateArea 2.600000 ;
    END I
    PIN OEN
        AntennaGateArea 2.730000 ;
    END OEN
    PIN PAD
        AntennaDiffArea 3461.000000 ;
    END PAD
END PRT12DGZ

MACRO PRT16DGZ
    PIN I
        AntennaGateArea 2.600000 ;
    END I
    PIN OEN
        AntennaGateArea 2.730000 ;
    END OEN
    PIN PAD
        AntennaDiffArea 3200.000000 ;
    END PAD
END PRT16DGZ

MACRO PDU02SDGZ
    PIN C
        AntennaDiffArea 3.660000 ;
    END C
    PIN I
        AntennaGateArea 2.600000 ;
    END I
    PIN OEN
        AntennaGateArea 2.730000 ;
    END OEN
    PIN PAD
        AntennaGateArea 4.800000 ;
        AntennaDiffArea 3670.000000 ;
    END PAD
END PDU02SDGZ

MACRO PRB08SDGZ
    PIN C
        AntennaDiffArea 3.660000 ;
    END C
    PIN I
        AntennaGateArea 2.600000 ;
    END I
    PIN OEN
        AntennaGateArea 2.730000 ;
    END OEN
    PIN PAD
        AntennaGateArea 4.800000 ;
        AntennaDiffArea 3486.000000 ;
    END PAD
END PRB08SDGZ

MACRO PRDW12DGZ
    PIN C
        AntennaDiffArea 3.660000 ;
    END C
    PIN I
        AntennaGateArea 2.600000 ;
    END I
    PIN OEN
        AntennaGateArea 2.730000 ;
    END OEN
    PIN PAD
        AntennaGateArea 3.600000 ;
        AntennaDiffArea 3478.000000 ;
    END PAD
    PIN REN
        AntennaGateArea 1.170000 ;
    END REN
END PRDW12DGZ

MACRO PDU04SDGZ
    PIN C
        AntennaDiffArea 3.660000 ;
    END C
    PIN I
        AntennaGateArea 2.600000 ;
    END I
    PIN OEN
        AntennaGateArea 2.730000 ;
    END OEN
    PIN PAD
        AntennaGateArea 4.800000 ;
        AntennaDiffArea 3484.000000 ;
    END PAD
END PDU04SDGZ

MACRO PRD08SDGZ
    PIN C
        AntennaDiffArea 3.660000 ;
    END C
    PIN I
        AntennaGateArea 2.600000 ;
    END I
    PIN OEN
        AntennaGateArea 2.730000 ;
    END OEN
    PIN PAD
        AntennaGateArea 4.800000 ;
        AntennaDiffArea 3486.000000 ;
    END PAD
END PRD08SDGZ

MACRO PDXO01DG
    PIN XC
        AntennaDiffArea 6.720000 ;
    END XC
    PIN XIN
        AntennaGateArea 220.000000 ;
        AntennaDiffArea 4126.000000 ;
    END XIN
    PIN XOUT
        AntennaGateArea 28.000000 ;
        AntennaDiffArea 2965.000000 ;
    END XOUT
END PDXO01DG

MACRO PDUW02DGZ
    PIN C
        AntennaDiffArea 3.660000 ;
    END C
    PIN I
        AntennaGateArea 2.600000 ;
    END I
    PIN OEN
        AntennaGateArea 2.730000 ;
    END OEN
    PIN PAD
        AntennaGateArea 3.600000 ;
        AntennaDiffArea 3670.000000 ;
    END PAD
    PIN REN
        AntennaGateArea 8.170000 ;
    END REN
END PDUW02DGZ

MACRO PDUW12DGZ
    PIN C
        AntennaDiffArea 3.660000 ;
    END C
    PIN I
        AntennaGateArea 2.600000 ;
    END I
    PIN OEN
        AntennaGateArea 2.730000 ;
    END OEN
    PIN PAD
        AntennaGateArea 3.600000 ;
        AntennaDiffArea 3478.000000 ;
    END PAD
    PIN REN
        AntennaGateArea 8.170000 ;
    END REN
END PDUW12DGZ

MACRO PRDW16DGZ
    PIN C
        AntennaDiffArea 3.660000 ;
    END C
    PIN I
        AntennaGateArea 2.600000 ;
    END I
    PIN OEN
        AntennaGateArea 2.730000 ;
    END OEN
    PIN PAD
        AntennaGateArea 3.600000 ;
        AntennaDiffArea 3217.000000 ;
    END PAD
    PIN REN
        AntennaGateArea 1.170000 ;
    END REN
END PRDW16DGZ

MACRO PDXO03DG
    PIN XC
        AntennaDiffArea 6.720000 ;
    END XC
    PIN XIN
        AntennaGateArea 205.000000 ;
        AntennaDiffArea 4126.000000 ;
    END XIN
    PIN XOUT
        AntennaGateArea 28.000000 ;
        AntennaDiffArea 3413.000000 ;
    END XOUT
END PDXO03DG

MACRO PDU08SDGZ
    PIN C
        AntennaDiffArea 3.660000 ;
    END C
    PIN I
        AntennaGateArea 2.600000 ;
    END I
    PIN OEN
        AntennaGateArea 2.730000 ;
    END OEN
    PIN PAD
        AntennaGateArea 4.800000 ;
        AntennaDiffArea 3486.000000 ;
    END PAD
END PDU08SDGZ

MACRO PDUW16DGZ
    PIN C
        AntennaDiffArea 3.660000 ;
    END C
    PIN I
        AntennaGateArea 2.600000 ;
    END I
    PIN OEN
        AntennaGateArea 2.730000 ;
    END OEN
    PIN PAD
        AntennaGateArea 3.600000 ;
        AntennaDiffArea 3217.000000 ;
    END PAD
    PIN REN
        AntennaGateArea 8.170000 ;
    END REN
END PDUW16DGZ

MACRO PDU02DGZ
    PIN C
        AntennaDiffArea 3.660000 ;
    END C
    PIN I
        AntennaGateArea 2.600000 ;
    END I
    PIN OEN
        AntennaGateArea 2.730000 ;
    END OEN
    PIN PAD
        AntennaGateArea 3.600000 ;
        AntennaDiffArea 3670.000000 ;
    END PAD
END PDU02DGZ

MACRO PDU12DGZ
    PIN C
        AntennaDiffArea 3.660000 ;
    END C
    PIN I
        AntennaGateArea 2.600000 ;
    END I
    PIN OEN
        AntennaGateArea 2.730000 ;
    END OEN
    PIN PAD
        AntennaGateArea 3.600000 ;
        AntennaDiffArea 3478.000000 ;
    END PAD
END PDU12DGZ

MACRO PDO02CDG
    PIN I
        AntennaGateArea 2.600000 ;
    END I
    PIN PAD
        AntennaDiffArea 4172.000000 ;
    END PAD
END PDO02CDG

MACRO PDO12CDG
    PIN I
        AntennaGateArea 2.600000 ;
    END I
    PIN PAD
        AntennaDiffArea 3963.000000 ;
    END PAD
END PDO12CDG

MACRO PRU24SDGZ
    PIN C
        AntennaDiffArea 3.660000 ;
    END C
    PIN I
        AntennaGateArea 2.600000 ;
    END I
    PIN OEN
        AntennaGateArea 2.730000 ;
    END OEN
    PIN PAD
        AntennaGateArea 4.800000 ;
        AntennaDiffArea 3479.000000 ;
    END PAD
END PRU24SDGZ

MACRO PDU16DGZ
    PIN C
        AntennaDiffArea 3.660000 ;
    END C
    PIN I
        AntennaGateArea 2.600000 ;
    END I
    PIN OEN
        AntennaGateArea 2.730000 ;
    END OEN
    PIN PAD
        AntennaGateArea 3.600000 ;
        AntennaDiffArea 3217.000000 ;
    END PAD
END PDU16DGZ

MACRO PDO16CDG
    PIN I
        AntennaGateArea 2.600000 ;
    END I
    PIN PAD
        AntennaDiffArea 3659.000000 ;
    END PAD
END PDO16CDG

MACRO PRUW24DGZ
    PIN C
        AntennaDiffArea 3.660000 ;
    END C
    PIN I
        AntennaGateArea 2.600000 ;
    END I
    PIN OEN
        AntennaGateArea 2.730000 ;
    END OEN
    PIN PAD
        AntennaGateArea 3.600000 ;
        AntennaDiffArea 3479.000000 ;
    END PAD
    PIN REN
        AntennaGateArea 8.170000 ;
    END REN
END PRUW24DGZ

MACRO PRUW08DGZ
    PIN C
        AntennaDiffArea 3.660000 ;
    END C
    PIN I
        AntennaGateArea 2.600000 ;
    END I
    PIN OEN
        AntennaGateArea 2.730000 ;
    END OEN
    PIN PAD
        AntennaGateArea 3.600000 ;
        AntennaDiffArea 3486.000000 ;
    END PAD
    PIN REN
        AntennaGateArea 8.170000 ;
    END REN
END PRUW08DGZ

MACRO PDXOE1DG
    PIN E
        AntennaGateArea 8.350000 ;
    END E
    PIN XC
        AntennaDiffArea 6.720000 ;
    END XC
    PIN XIN
        AntennaGateArea 200.000000 ;
        AntennaDiffArea 4126.000000 ;
    END XIN
    PIN XOUT
        AntennaGateArea 28.000000 ;
        AntennaDiffArea 2968.000000 ;
    END XOUT
END PDXOE1DG

MACRO PDB02DGZ
    PIN C
        AntennaDiffArea 3.660000 ;
    END C
    PIN I
        AntennaGateArea 2.600000 ;
    END I
    PIN OEN
        AntennaGateArea 2.730000 ;
    END OEN
    PIN PAD
        AntennaGateArea 3.600000 ;
        AntennaDiffArea 3670.000000 ;
    END PAD
END PDB02DGZ

MACRO PDXOE3DG
    PIN E
        AntennaGateArea 8.350000 ;
    END E
    PIN XC
        AntennaDiffArea 6.720000 ;
    END XC
    PIN XIN
        AntennaGateArea 125.000000 ;
        AntennaDiffArea 4126.000000 ;
    END XIN
    PIN XOUT
        AntennaGateArea 28.000000 ;
        AntennaDiffArea 3638.000000 ;
    END XOUT
END PDXOE3DG

MACRO PDB12DGZ
    PIN C
        AntennaDiffArea 3.660000 ;
    END C
    PIN I
        AntennaGateArea 2.600000 ;
    END I
    PIN OEN
        AntennaGateArea 2.730000 ;
    END OEN
    PIN PAD
        AntennaGateArea 3.600000 ;
        AntennaDiffArea 3478.000000 ;
    END PAD
END PDB12DGZ

MACRO PRU12DGZ
    PIN C
        AntennaDiffArea 3.660000 ;
    END C
    PIN I
        AntennaGateArea 2.600000 ;
    END I
    PIN OEN
        AntennaGateArea 2.730000 ;
    END OEN
    PIN PAD
        AntennaGateArea 3.600000 ;
        AntennaDiffArea 3478.000000 ;
    END PAD
END PRU12DGZ

MACRO PRB12SDGZ
    PIN C
        AntennaDiffArea 3.660000 ;
    END C
    PIN I
        AntennaGateArea 2.600000 ;
    END I
    PIN OEN
        AntennaGateArea 2.730000 ;
    END OEN
    PIN PAD
        AntennaGateArea 4.800000 ;
        AntennaDiffArea 3478.000000 ;
    END PAD
END PRB12SDGZ

MACRO PRD12SDGZ
    PIN C
        AntennaDiffArea 3.660000 ;
    END C
    PIN I
        AntennaGateArea 2.600000 ;
    END I
    PIN OEN
        AntennaGateArea 2.730000 ;
    END OEN
    PIN PAD
        AntennaGateArea 4.800000 ;
        AntennaDiffArea 3478.000000 ;
    END PAD
END PRD12SDGZ

MACRO PDD04DGZ
    PIN C
        AntennaDiffArea 3.660000 ;
    END C
    PIN I
        AntennaGateArea 2.600000 ;
    END I
    PIN OEN
        AntennaGateArea 2.730000 ;
    END OEN
    PIN PAD
        AntennaGateArea 3.600000 ;
        AntennaDiffArea 3484.000000 ;
    END PAD
END PDD04DGZ

MACRO PRO12CDG
    PIN I
        AntennaGateArea 2.600000 ;
    END I
    PIN PAD
        AntennaDiffArea 3963.000000 ;
    END PAD
END PRO12CDG

MACRO PDB16DGZ
    PIN C
        AntennaDiffArea 3.660000 ;
    END C
    PIN I
        AntennaGateArea 2.600000 ;
    END I
    PIN OEN
        AntennaGateArea 2.730000 ;
    END OEN
    PIN PAD
        AntennaGateArea 3.600000 ;
        AntennaDiffArea 3217.000000 ;
    END PAD
END PDB16DGZ

MACRO PDIDGZ
    PIN C
        AntennaDiffArea 3.660000 ;
    END C
    PIN PAD
        AntennaGateArea 3.600000 ;
        AntennaDiffArea 3670.000000 ;
    END PAD
END PDIDGZ

MACRO PRU16DGZ
    PIN C
        AntennaDiffArea 3.660000 ;
    END C
    PIN I
        AntennaGateArea 2.600000 ;
    END I
    PIN OEN
        AntennaGateArea 2.730000 ;
    END OEN
    PIN PAD
        AntennaGateArea 3.600000 ;
        AntennaDiffArea 3217.000000 ;
    END PAD
END PRU16DGZ

MACRO PRB16SDGZ
    PIN C
        AntennaDiffArea 3.660000 ;
    END C
    PIN I
        AntennaGateArea 2.600000 ;
    END I
    PIN OEN
        AntennaGateArea 2.730000 ;
    END OEN
    PIN PAD
        AntennaGateArea 4.800000 ;
        AntennaDiffArea 3217.000000 ;
    END PAD
END PRB16SDGZ

MACRO PDD24DGZ
    PIN C
        AntennaDiffArea 3.660000 ;
    END C
    PIN I
        AntennaGateArea 2.600000 ;
    END I
    PIN OEN
        AntennaGateArea 2.730000 ;
    END OEN
    PIN PAD
        AntennaGateArea 3.600000 ;
        AntennaDiffArea 3479.000000 ;
    END PAD
END PDD24DGZ

MACRO PDU12SDGZ
    PIN C
        AntennaDiffArea 3.660000 ;
    END C
    PIN I
        AntennaGateArea 2.600000 ;
    END I
    PIN OEN
        AntennaGateArea 2.730000 ;
    END OEN
    PIN PAD
        AntennaGateArea 4.800000 ;
        AntennaDiffArea 3478.000000 ;
    END PAD
END PDU12SDGZ

MACRO PRD16SDGZ
    PIN C
        AntennaDiffArea 3.660000 ;
    END C
    PIN I
        AntennaGateArea 2.600000 ;
    END I
    PIN OEN
        AntennaGateArea 2.730000 ;
    END OEN
    PIN PAD
        AntennaGateArea 4.800000 ;
        AntennaDiffArea 3217.000000 ;
    END PAD
END PRD16SDGZ

MACRO PDD08DGZ
    PIN C
        AntennaDiffArea 3.660000 ;
    END C
    PIN I
        AntennaGateArea 2.600000 ;
    END I
    PIN OEN
        AntennaGateArea 2.730000 ;
    END OEN
    PIN PAD
        AntennaGateArea 3.600000 ;
        AntennaDiffArea 3486.000000 ;
    END PAD
END PDD08DGZ

MACRO PRO16CDG
    PIN I
        AntennaGateArea 2.600000 ;
    END I
    PIN PAD
        AntennaDiffArea 3659.000000 ;
    END PAD
END PRO16CDG

MACRO PDU16SDGZ
    PIN C
        AntennaDiffArea 3.660000 ;
    END C
    PIN I
        AntennaGateArea 2.600000 ;
    END I
    PIN OEN
        AntennaGateArea 2.730000 ;
    END OEN
    PIN PAD
        AntennaGateArea 4.800000 ;
        AntennaDiffArea 3217.000000 ;
    END PAD
END PDU16SDGZ

MACRO PRB12DGZ
    PIN C
        AntennaDiffArea 3.660000 ;
    END C
    PIN I
        AntennaGateArea 2.600000 ;
    END I
    PIN OEN
        AntennaGateArea 2.730000 ;
    END OEN
    PIN PAD
        AntennaGateArea 3.600000 ;
        AntennaDiffArea 3478.000000 ;
    END PAD
END PRB12DGZ

MACRO PDUDGZ
    PIN C
        AntennaDiffArea 3.660000 ;
    END C
    PIN PAD
        AntennaGateArea 3.600000 ;
        AntennaDiffArea 3670.000000 ;
    END PAD
END PDUDGZ

MACRO PRB16DGZ
    PIN C
        AntennaDiffArea 3.660000 ;
    END C
    PIN I
        AntennaGateArea 2.600000 ;
    END I
    PIN OEN
        AntennaGateArea 2.730000 ;
    END OEN
    PIN PAD
        AntennaGateArea 3.600000 ;
        AntennaDiffArea 3217.000000 ;
    END PAD
END PRB16DGZ

MACRO PDB02SDGZ
    PIN C
        AntennaDiffArea 3.660000 ;
    END C
    PIN I
        AntennaGateArea 2.600000 ;
    END I
    PIN OEN
        AntennaGateArea 2.730000 ;
    END OEN
    PIN PAD
        AntennaGateArea 4.800000 ;
        AntennaDiffArea 3670.000000 ;
    END PAD
END PDB02SDGZ

MACRO PRD24DGZ
    PIN C
        AntennaDiffArea 3.660000 ;
    END C
    PIN I
        AntennaGateArea 2.600000 ;
    END I
    PIN OEN
        AntennaGateArea 2.730000 ;
    END OEN
    PIN PAD
        AntennaGateArea 3.600000 ;
        AntennaDiffArea 3479.000000 ;
    END PAD
END PRD24DGZ

MACRO PDT04DGZ
    PIN I
        AntennaGateArea 2.600000 ;
    END I
    PIN OEN
        AntennaGateArea 2.730000 ;
    END OEN
    PIN PAD
        AntennaDiffArea 3467.000000 ;
    END PAD
END PDT04DGZ

MACRO PDD02SDGZ
    PIN C
        AntennaDiffArea 3.660000 ;
    END C
    PIN I
        AntennaGateArea 2.600000 ;
    END I
    PIN OEN
        AntennaGateArea 2.730000 ;
    END OEN
    PIN PAD
        AntennaGateArea 4.800000 ;
        AntennaDiffArea 3670.000000 ;
    END PAD
END PDD02SDGZ

MACRO PDB04SDGZ
    PIN C
        AntennaDiffArea 3.660000 ;
    END C
    PIN I
        AntennaGateArea 2.600000 ;
    END I
    PIN OEN
        AntennaGateArea 2.730000 ;
    END OEN
    PIN PAD
        AntennaGateArea 4.800000 ;
        AntennaDiffArea 3484.000000 ;
    END PAD
END PDB04SDGZ

MACRO PRD08DGZ
    PIN C
        AntennaDiffArea 3.660000 ;
    END C
    PIN I
        AntennaGateArea 2.600000 ;
    END I
    PIN OEN
        AntennaGateArea 2.730000 ;
    END OEN
    PIN PAD
        AntennaGateArea 3.600000 ;
        AntennaDiffArea 3486.000000 ;
    END PAD
END PRD08DGZ

MACRO PDT24DGZ
    PIN I
        AntennaGateArea 2.600000 ;
    END I
    PIN OEN
        AntennaGateArea 2.730000 ;
    END OEN
    PIN PAD
        AntennaDiffArea 3461.000000 ;
    END PAD
END PDT24DGZ

MACRO PDD04SDGZ
    PIN C
        AntennaDiffArea 3.660000 ;
    END C
    PIN I
        AntennaGateArea 2.600000 ;
    END I
    PIN OEN
        AntennaGateArea 2.730000 ;
    END OEN
    PIN PAD
        AntennaGateArea 4.800000 ;
        AntennaDiffArea 3484.000000 ;
    END PAD
END PDD04SDGZ

MACRO PDT08DGZ
    PIN I
        AntennaGateArea 2.600000 ;
    END I
    PIN OEN
        AntennaGateArea 2.730000 ;
    END OEN
    PIN PAD
        AntennaDiffArea 3469.000000 ;
    END PAD
END PDT08DGZ

MACRO PDB08SDGZ
    PIN C
        AntennaDiffArea 3.660000 ;
    END C
    PIN I
        AntennaGateArea 2.600000 ;
    END I
    PIN OEN
        AntennaGateArea 2.730000 ;
    END OEN
    PIN PAD
        AntennaGateArea 4.800000 ;
        AntennaDiffArea 3486.000000 ;
    END PAD
END PDB08SDGZ

MACRO PDDW02DGZ
    PIN C
        AntennaDiffArea 3.660000 ;
    END C
    PIN I
        AntennaGateArea 2.600000 ;
    END I
    PIN OEN
        AntennaGateArea 2.730000 ;
    END OEN
    PIN PAD
        AntennaGateArea 3.600000 ;
        AntennaDiffArea 3670.000000 ;
    END PAD
    PIN REN
        AntennaGateArea 1.170000 ;
    END REN
END PDDW02DGZ

MACRO PDDW12DGZ
    PIN C
        AntennaDiffArea 3.660000 ;
    END C
    PIN I
        AntennaGateArea 2.600000 ;
    END I
    PIN OEN
        AntennaGateArea 2.730000 ;
    END OEN
    PIN PAD
        AntennaGateArea 3.600000 ;
        AntennaDiffArea 3478.000000 ;
    END PAD
    PIN REN
        AntennaGateArea 1.170000 ;
    END REN
END PDDW12DGZ

MACRO PDD08SDGZ
    PIN C
        AntennaDiffArea 3.660000 ;
    END C
    PIN I
        AntennaGateArea 2.600000 ;
    END I
    PIN OEN
        AntennaGateArea 2.730000 ;
    END OEN
    PIN PAD
        AntennaGateArea 4.800000 ;
        AntennaDiffArea 3486.000000 ;
    END PAD
END PDD08SDGZ

MACRO PDDW16DGZ
    PIN C
        AntennaDiffArea 3.660000 ;
    END C
    PIN I
        AntennaGateArea 2.600000 ;
    END I
    PIN OEN
        AntennaGateArea 2.730000 ;
    END OEN
    PIN PAD
        AntennaGateArea 3.600000 ;
        AntennaDiffArea 3217.000000 ;
    END PAD
    PIN REN
        AntennaGateArea 1.170000 ;
    END REN
END PDDW16DGZ

MACRO PDDDGZ
    PIN C
        AntennaDiffArea 3.660000 ;
    END C
    PIN PAD
        AntennaGateArea 3.600000 ;
        AntennaDiffArea 3670.000000 ;
    END PAD
END PDDDGZ

MACRO PRT24DGZ
    PIN I
        AntennaGateArea 2.600000 ;
    END I
    PIN OEN
        AntennaGateArea 2.730000 ;
    END OEN
    PIN PAD
        AntennaDiffArea 3461.000000 ;
    END PAD
END PRT24DGZ

MACRO PVSS1DGZ
    PIN VSS
        AntennaDiffArea 1996.000000 ;
    END VSS
END PVSS1DGZ

MACRO PRB24SDGZ
    PIN C
        AntennaDiffArea 3.660000 ;
    END C
    PIN I
        AntennaGateArea 2.600000 ;
    END I
    PIN OEN
        AntennaGateArea 2.730000 ;
    END OEN
    PIN PAD
        AntennaGateArea 4.800000 ;
        AntennaDiffArea 3479.000000 ;
    END PAD
END PRB24SDGZ

MACRO PRT08DGZ
    PIN I
        AntennaGateArea 2.600000 ;
    END I
    PIN OEN
        AntennaGateArea 2.730000 ;
    END OEN
    PIN PAD
        AntennaDiffArea 3469.000000 ;
    END PAD
END PRT08DGZ

MACRO PVDD1DGZ
    PIN VDD
        AntennaDiffArea 4389.000000 ;
    END VDD
END PVDD1DGZ

MACRO PRD24SDGZ
    PIN C
        AntennaDiffArea 3.660000 ;
    END C
    PIN I
        AntennaGateArea 2.600000 ;
    END I
    PIN OEN
        AntennaGateArea 2.730000 ;
    END OEN
    PIN PAD
        AntennaGateArea 4.800000 ;
        AntennaDiffArea 3479.000000 ;
    END PAD
END PRD24SDGZ

MACRO PDU24SDGZ
    PIN C
        AntennaDiffArea 3.660000 ;
    END C
    PIN I
        AntennaGateArea 2.600000 ;
    END I
    PIN OEN
        AntennaGateArea 2.730000 ;
    END OEN
    PIN PAD
        AntennaGateArea 4.800000 ;
        AntennaDiffArea 3479.000000 ;
    END PAD
END PDU24SDGZ

MACRO PRDW24DGZ
    PIN C
        AntennaDiffArea 3.660000 ;
    END C
    PIN I
        AntennaGateArea 2.600000 ;
    END I
    PIN OEN
        AntennaGateArea 2.730000 ;
    END OEN
    PIN PAD
        AntennaGateArea 3.600000 ;
        AntennaDiffArea 3479.000000 ;
    END PAD
    PIN REN
        AntennaGateArea 1.170000 ;
    END REN
END PRDW24DGZ

MACRO PDXO02DG
    PIN XC
        AntennaDiffArea 6.720000 ;
    END XC
    PIN XIN
        AntennaGateArea 170.000000 ;
        AntennaDiffArea 4126.000000 ;
    END XIN
    PIN XOUT
        AntennaGateArea 28.000000 ;
        AntennaDiffArea 3101.000000 ;
    END XOUT
END PDXO02DG

MACRO PDUW04DGZ
    PIN C
        AntennaDiffArea 3.660000 ;
    END C
    PIN I
        AntennaGateArea 2.600000 ;
    END I
    PIN OEN
        AntennaGateArea 2.730000 ;
    END OEN
    PIN PAD
        AntennaGateArea 3.600000 ;
        AntennaDiffArea 3484.000000 ;
    END PAD
    PIN REN
        AntennaGateArea 8.170000 ;
    END REN
END PDUW04DGZ

MACRO PRDW08DGZ
    PIN C
        AntennaDiffArea 3.660000 ;
    END C
    PIN I
        AntennaGateArea 2.600000 ;
    END I
    PIN OEN
        AntennaGateArea 2.730000 ;
    END OEN
    PIN PAD
        AntennaGateArea 3.600000 ;
        AntennaDiffArea 3486.000000 ;
    END PAD
    PIN REN
        AntennaGateArea 1.170000 ;
    END REN
END PRDW08DGZ

MACRO PDUW24DGZ
    PIN C
        AntennaDiffArea 3.660000 ;
    END C
    PIN I
        AntennaGateArea 2.600000 ;
    END I
    PIN OEN
        AntennaGateArea 2.730000 ;
    END OEN
    PIN PAD
        AntennaGateArea 3.600000 ;
        AntennaDiffArea 3479.000000 ;
    END PAD
    PIN REN
        AntennaGateArea 8.170000 ;
    END REN
END PDUW24DGZ

MACRO PDUW08DGZ
    PIN C
        AntennaDiffArea 3.660000 ;
    END C
    PIN I
        AntennaGateArea 2.600000 ;
    END I
    PIN OEN
        AntennaGateArea 2.730000 ;
    END OEN
    PIN PAD
        AntennaGateArea 3.600000 ;
        AntennaDiffArea 3486.000000 ;
    END PAD
    PIN REN
        AntennaGateArea 8.170000 ;
    END REN
END PDUW08DGZ

MACRO PDDSDGZ
    PIN C
        AntennaDiffArea 3.660000 ;
    END C
    PIN PAD
        AntennaGateArea 4.800000 ;
        AntennaDiffArea 3670.000000 ;
    END PAD
END PDDSDGZ

MACRO PDB12SDGZ
    PIN C
        AntennaDiffArea 3.660000 ;
    END C
    PIN I
        AntennaGateArea 2.600000 ;
    END I
    PIN OEN
        AntennaGateArea 2.730000 ;
    END OEN
    PIN PAD
        AntennaGateArea 4.800000 ;
        AntennaDiffArea 3478.000000 ;
    END PAD
END PDB12SDGZ

MACRO PDU04DGZ
    PIN C
        AntennaDiffArea 3.660000 ;
    END C
    PIN I
        AntennaGateArea 2.600000 ;
    END I
    PIN OEN
        AntennaGateArea 2.730000 ;
    END OEN
    PIN PAD
        AntennaGateArea 3.600000 ;
        AntennaDiffArea 3484.000000 ;
    END PAD
END PDU04DGZ

MACRO PDD12SDGZ
    PIN C
        AntennaDiffArea 3.660000 ;
    END C
    PIN I
        AntennaGateArea 2.600000 ;
    END I
    PIN OEN
        AntennaGateArea 2.730000 ;
    END OEN
    PIN PAD
        AntennaGateArea 4.800000 ;
        AntennaDiffArea 3478.000000 ;
    END PAD
END PDD12SDGZ

MACRO PDDWDGZ
    PIN C
        AntennaDiffArea 3.660000 ;
    END C
    PIN PAD
        AntennaGateArea 3.600000 ;
        AntennaDiffArea 3670.000000 ;
    END PAD
    PIN REN
        AntennaGateArea 1.170000 ;
    END REN
END PDDWDGZ

MACRO PDU24DGZ
    PIN C
        AntennaDiffArea 3.660000 ;
    END C
    PIN I
        AntennaGateArea 2.600000 ;
    END I
    PIN OEN
        AntennaGateArea 2.730000 ;
    END OEN
    PIN PAD
        AntennaGateArea 3.600000 ;
        AntennaDiffArea 3479.000000 ;
    END PAD
END PDU24DGZ

MACRO PDB16SDGZ
    PIN C
        AntennaDiffArea 3.660000 ;
    END C
    PIN I
        AntennaGateArea 2.600000 ;
    END I
    PIN OEN
        AntennaGateArea 2.730000 ;
    END OEN
    PIN PAD
        AntennaGateArea 4.800000 ;
        AntennaDiffArea 3217.000000 ;
    END PAD
END PDB16SDGZ

MACRO PDISDGZ
    PIN C
        AntennaDiffArea 3.660000 ;
    END C
    PIN PAD
        AntennaGateArea 4.800000 ;
        AntennaDiffArea 3670.000000 ;
    END PAD
END PDISDGZ

MACRO PDO04CDG
    PIN I
        AntennaGateArea 2.600000 ;
    END I
    PIN PAD
        AntennaDiffArea 4072.000000 ;
    END PAD
END PDO04CDG

MACRO PRUW12DGZ
    PIN C
        AntennaDiffArea 3.660000 ;
    END C
    PIN I
        AntennaGateArea 2.600000 ;
    END I
    PIN OEN
        AntennaGateArea 2.730000 ;
    END OEN
    PIN PAD
        AntennaGateArea 3.600000 ;
        AntennaDiffArea 3478.000000 ;
    END PAD
    PIN REN
        AntennaGateArea 8.170000 ;
    END REN
END PRUW12DGZ

MACRO PDU08DGZ
    PIN C
        AntennaDiffArea 3.660000 ;
    END C
    PIN I
        AntennaGateArea 2.600000 ;
    END I
    PIN OEN
        AntennaGateArea 2.730000 ;
    END OEN
    PIN PAD
        AntennaGateArea 3.600000 ;
        AntennaDiffArea 3486.000000 ;
    END PAD
END PDU08DGZ

MACRO PRU08SDGZ
    PIN C
        AntennaDiffArea 3.660000 ;
    END C
    PIN I
        AntennaGateArea 2.600000 ;
    END I
    PIN OEN
        AntennaGateArea 2.730000 ;
    END OEN
    PIN PAD
        AntennaGateArea 4.800000 ;
        AntennaDiffArea 3486.000000 ;
    END PAD
END PRU08SDGZ

MACRO PDD16SDGZ
    PIN C
        AntennaDiffArea 3.660000 ;
    END C
    PIN I
        AntennaGateArea 2.600000 ;
    END I
    PIN OEN
        AntennaGateArea 2.730000 ;
    END OEN
    PIN PAD
        AntennaGateArea 4.800000 ;
        AntennaDiffArea 3217.000000 ;
    END PAD
END PDD16SDGZ

MACRO PDO24CDG
    PIN I
        AntennaGateArea 2.600000 ;
    END I
    PIN PAD
        AntennaDiffArea 4047.000000 ;
    END PAD
END PDO24CDG

MACRO PDO08CDG
    PIN I
        AntennaGateArea 2.600000 ;
    END I
    PIN PAD
        AntennaDiffArea 4037.000000 ;
    END PAD
END PDO08CDG

MACRO PRUW16DGZ
    PIN C
        AntennaDiffArea 3.660000 ;
    END C
    PIN I
        AntennaGateArea 2.600000 ;
    END I
    PIN OEN
        AntennaGateArea 2.730000 ;
    END OEN
    PIN PAD
        AntennaGateArea 3.600000 ;
        AntennaDiffArea 3217.000000 ;
    END PAD
    PIN REN
        AntennaGateArea 8.170000 ;
    END REN
END PRUW16DGZ

MACRO PDXOE2DG
    PIN E
        AntennaGateArea 8.350000 ;
    END E
    PIN XC
        AntennaDiffArea 6.720000 ;
    END XC
    PIN XIN
        AntennaGateArea 130.000000 ;
        AntennaDiffArea 4126.000000 ;
    END XIN
    PIN XOUT
        AntennaGateArea 28.000000 ;
        AntennaDiffArea 3278.000000 ;
    END XOUT
END PDXOE2DG

MACRO PDB04DGZ
    PIN C
        AntennaDiffArea 3.660000 ;
    END C
    PIN I
        AntennaGateArea 2.600000 ;
    END I
    PIN OEN
        AntennaGateArea 2.730000 ;
    END OEN
    PIN PAD
        AntennaGateArea 3.600000 ;
        AntennaDiffArea 3484.000000 ;
    END PAD
END PDB04DGZ

MACRO PDD02DGZ
    PIN C
        AntennaDiffArea 3.660000 ;
    END C
    PIN I
        AntennaGateArea 2.600000 ;
    END I
    PIN OEN
        AntennaGateArea 2.730000 ;
    END OEN
    PIN PAD
        AntennaGateArea 3.600000 ;
        AntennaDiffArea 3670.000000 ;
    END PAD
END PDD02DGZ

END LIBRARY
